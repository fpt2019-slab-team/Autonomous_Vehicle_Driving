//-----------------------------------------------------------------------------
// <arctan_calc> 
//  - Pipelined arctangent calculation module
//    - behaves like numpy.arctan2(in_x1, in_x2)
//    - <in_x1>, <in_x2>: 9-bit signed coordinates
//    - <out_val>: [0, 256) (equivalent to [0, 2pi))
//  - Overall latency is 5 clock cycles
//-----------------------------------------------------------------------------
// Version 1.00 (Oct. 30, 2019)
//  - Initial version
//-----------------------------------------------------------------------------
// (C) 2019 Taito Manabe. All rights reserved.
//-----------------------------------------------------------------------------
`default_nettype none
`timescale 1ns/1ns
  
module arctan_calc
  ( clock, in_x1, in_x2, out_val );

   // inputs/outputs ----------------------------------------------------------
   input wire       	   clock;
   input wire signed [8:0] in_x1, in_x2;
   output reg [7:0] 	   out_val;

   // -------------------------------------------------------------------------
   // [stage 1] condition check
   reg 	      s1_x_zero, s1_y_zero, s1_x_neg, s1_y_neg;
   reg [7:0]  s1_x, s1_y;
   always @(posedge clock) begin
      s1_x <= absolute(in_x1);
      s1_y <= absolute(in_x2);
      s1_x_zero <= (in_x1 == 0);
      s1_y_zero <= (in_x2 == 0);
      s1_x_neg  <= (in_x1  < 0);
      s1_y_neg  <= (in_x2  < 0);
   end

   // [stage 2] preparation for address calculation
   reg        s2_x_zero, s2_y_zero, s2_x_neg, s2_y_neg, s2_swap;
   reg [5:0]  s2_x, s2_y;
   always @(posedge clock) begin
      {s2_x_zero, s2_y_zero, s2_x_neg, s2_y_neg}
	<= {s1_x_zero, s1_y_zero, s1_x_neg, s1_y_neg};
      if(s1_y < s1_x) begin
	 s2_swap <= 1;
	 if(s1_x < 64)
	   {s2_x, s2_y} <= {s1_y[5:0], s1_x[5:0]};
	 else if(s1_x < 128)
	   {s2_x, s2_y} <= {s1_y[6:1], s1_x[6:1]};
	 else
	   {s2_x, s2_y} <= {s1_y[7:2], s1_x[7:2]};
      end
      else begin
	 s2_swap <= 0;
	 if(s1_y < 64)
	   {s2_x, s2_y} <= {s1_x[5:0], s1_y[5:0]};
	 else if(s1_y < 128)
	   {s2_x, s2_y} <= {s1_x[6:1], s1_y[6:1]};
	 else
	   {s2_x, s2_y} <= {s1_x[7:2], s1_y[7:2]};
      end
   end

   // [stage 3] address calculation
   reg        s3_x_zero, s3_y_zero, s3_x_neg, s3_y_neg, s3_swap, s3_match;
   reg [10:0] s3_addr;
   always @(posedge clock) begin
      {s3_x_zero, s3_y_zero, s3_x_neg, s3_y_neg, s3_swap}
	<= {s2_x_zero, s2_y_zero, s2_x_neg, s2_y_neg, s2_swap};
      s3_match <= (s2_x == s2_y);
      if(s2_x_zero || s2_y_zero)
	s3_addr <= 0;  // don't care
      else
	s3_addr <= s2_y * (s2_y - 1) / 2 + s2_x - 1;
   end

   // [stage 4] reads data from ROM
   reg        s4_x_zero, s4_y_zero, s4_x_neg, s4_y_neg, s4_swap, s4_match;
   reg [4:0]  s4_angle;
   always @(posedge clock) begin
      {s4_x_zero, s4_y_zero, s4_x_neg, s4_y_neg, s4_swap, s4_match}
	<= {s3_x_zero, s3_y_zero, s3_x_neg, s3_y_neg, s3_swap, s3_match};
      case(s3_addr)
        0: s4_angle <= 0;
        1: s4_angle <= 19;
        2: s4_angle <= 0;
        3: s4_angle <= 13;
        4: s4_angle <= 24;
        5: s4_angle <= 0;
        6: s4_angle <= 10;
        7: s4_angle <= 19;
        8: s4_angle <= 26;
        9: s4_angle <= 0;
        10: s4_angle <= 8;
        11: s4_angle <= 16;
        12: s4_angle <= 22;
        13: s4_angle <= 27;
        14: s4_angle <= 0;
        15: s4_angle <= 7;
        16: s4_angle <= 13;
        17: s4_angle <= 19;
        18: s4_angle <= 24;
        19: s4_angle <= 28;
        20: s4_angle <= 0;
        21: s4_angle <= 6;
        22: s4_angle <= 11;
        23: s4_angle <= 16;
        24: s4_angle <= 21;
        25: s4_angle <= 25;
        26: s4_angle <= 29;
        27: s4_angle <= 0;
        28: s4_angle <= 5;
        29: s4_angle <= 10;
        30: s4_angle <= 15;
        31: s4_angle <= 19;
        32: s4_angle <= 23;
        33: s4_angle <= 26;
        34: s4_angle <= 29;
        35: s4_angle <= 0;
        36: s4_angle <= 5;
        37: s4_angle <= 9;
        38: s4_angle <= 13;
        39: s4_angle <= 17;
        40: s4_angle <= 21;
        41: s4_angle <= 24;
        42: s4_angle <= 27;
        43: s4_angle <= 30;
        44: s4_angle <= 0;
        45: s4_angle <= 4;
        46: s4_angle <= 8;
        47: s4_angle <= 12;
        48: s4_angle <= 16;
        49: s4_angle <= 19;
        50: s4_angle <= 22;
        51: s4_angle <= 25;
        52: s4_angle <= 27;
        53: s4_angle <= 30;
        54: s4_angle <= 0;
        55: s4_angle <= 4;
        56: s4_angle <= 7;
        57: s4_angle <= 11;
        58: s4_angle <= 14;
        59: s4_angle <= 17;
        60: s4_angle <= 20;
        61: s4_angle <= 23;
        62: s4_angle <= 26;
        63: s4_angle <= 28;
        64: s4_angle <= 30;
        65: s4_angle <= 0;
        66: s4_angle <= 3;
        67: s4_angle <= 7;
        68: s4_angle <= 10;
        69: s4_angle <= 13;
        70: s4_angle <= 16;
        71: s4_angle <= 19;
        72: s4_angle <= 22;
        73: s4_angle <= 24;
        74: s4_angle <= 26;
        75: s4_angle <= 28;
        76: s4_angle <= 30;
        77: s4_angle <= 0;
        78: s4_angle <= 3;
        79: s4_angle <= 6;
        80: s4_angle <= 9;
        81: s4_angle <= 12;
        82: s4_angle <= 15;
        83: s4_angle <= 18;
        84: s4_angle <= 20;
        85: s4_angle <= 22;
        86: s4_angle <= 25;
        87: s4_angle <= 27;
        88: s4_angle <= 29;
        89: s4_angle <= 30;
        90: s4_angle <= 0;
        91: s4_angle <= 3;
        92: s4_angle <= 6;
        93: s4_angle <= 9;
        94: s4_angle <= 11;
        95: s4_angle <= 14;
        96: s4_angle <= 16;
        97: s4_angle <= 19;
        98: s4_angle <= 21;
        99: s4_angle <= 23;
        100: s4_angle <= 25;
        101: s4_angle <= 27;
        102: s4_angle <= 29;
        103: s4_angle <= 30;
        104: s4_angle <= 0;
        105: s4_angle <= 3;
        106: s4_angle <= 5;
        107: s4_angle <= 8;
        108: s4_angle <= 11;
        109: s4_angle <= 13;
        110: s4_angle <= 16;
        111: s4_angle <= 18;
        112: s4_angle <= 20;
        113: s4_angle <= 22;
        114: s4_angle <= 24;
        115: s4_angle <= 26;
        116: s4_angle <= 27;
        117: s4_angle <= 29;
        118: s4_angle <= 31;
        119: s4_angle <= 0;
        120: s4_angle <= 3;
        121: s4_angle <= 5;
        122: s4_angle <= 8;
        123: s4_angle <= 10;
        124: s4_angle <= 12;
        125: s4_angle <= 15;
        126: s4_angle <= 17;
        127: s4_angle <= 19;
        128: s4_angle <= 21;
        129: s4_angle <= 23;
        130: s4_angle <= 25;
        131: s4_angle <= 26;
        132: s4_angle <= 28;
        133: s4_angle <= 29;
        134: s4_angle <= 31;
        135: s4_angle <= 0;
        136: s4_angle <= 2;
        137: s4_angle <= 5;
        138: s4_angle <= 7;
        139: s4_angle <= 9;
        140: s4_angle <= 12;
        141: s4_angle <= 14;
        142: s4_angle <= 16;
        143: s4_angle <= 18;
        144: s4_angle <= 20;
        145: s4_angle <= 22;
        146: s4_angle <= 23;
        147: s4_angle <= 25;
        148: s4_angle <= 27;
        149: s4_angle <= 28;
        150: s4_angle <= 29;
        151: s4_angle <= 31;
        152: s4_angle <= 0;
        153: s4_angle <= 2;
        154: s4_angle <= 5;
        155: s4_angle <= 7;
        156: s4_angle <= 9;
        157: s4_angle <= 11;
        158: s4_angle <= 13;
        159: s4_angle <= 15;
        160: s4_angle <= 17;
        161: s4_angle <= 19;
        162: s4_angle <= 21;
        163: s4_angle <= 22;
        164: s4_angle <= 24;
        165: s4_angle <= 25;
        166: s4_angle <= 27;
        167: s4_angle <= 28;
        168: s4_angle <= 30;
        169: s4_angle <= 31;
        170: s4_angle <= 0;
        171: s4_angle <= 2;
        172: s4_angle <= 4;
        173: s4_angle <= 6;
        174: s4_angle <= 8;
        175: s4_angle <= 10;
        176: s4_angle <= 12;
        177: s4_angle <= 14;
        178: s4_angle <= 16;
        179: s4_angle <= 18;
        180: s4_angle <= 20;
        181: s4_angle <= 21;
        182: s4_angle <= 23;
        183: s4_angle <= 24;
        184: s4_angle <= 26;
        185: s4_angle <= 27;
        186: s4_angle <= 29;
        187: s4_angle <= 30;
        188: s4_angle <= 31;
        189: s4_angle <= 0;
        190: s4_angle <= 2;
        191: s4_angle <= 4;
        192: s4_angle <= 6;
        193: s4_angle <= 8;
        194: s4_angle <= 10;
        195: s4_angle <= 12;
        196: s4_angle <= 14;
        197: s4_angle <= 16;
        198: s4_angle <= 17;
        199: s4_angle <= 19;
        200: s4_angle <= 20;
        201: s4_angle <= 22;
        202: s4_angle <= 23;
        203: s4_angle <= 25;
        204: s4_angle <= 26;
        205: s4_angle <= 27;
        206: s4_angle <= 29;
        207: s4_angle <= 30;
        208: s4_angle <= 31;
        209: s4_angle <= 0;
        210: s4_angle <= 2;
        211: s4_angle <= 4;
        212: s4_angle <= 6;
        213: s4_angle <= 8;
        214: s4_angle <= 10;
        215: s4_angle <= 11;
        216: s4_angle <= 13;
        217: s4_angle <= 15;
        218: s4_angle <= 16;
        219: s4_angle <= 18;
        220: s4_angle <= 20;
        221: s4_angle <= 21;
        222: s4_angle <= 23;
        223: s4_angle <= 24;
        224: s4_angle <= 25;
        225: s4_angle <= 27;
        226: s4_angle <= 28;
        227: s4_angle <= 29;
        228: s4_angle <= 30;
        229: s4_angle <= 31;
        230: s4_angle <= 0;
        231: s4_angle <= 2;
        232: s4_angle <= 4;
        233: s4_angle <= 6;
        234: s4_angle <= 7;
        235: s4_angle <= 9;
        236: s4_angle <= 11;
        237: s4_angle <= 13;
        238: s4_angle <= 14;
        239: s4_angle <= 16;
        240: s4_angle <= 17;
        241: s4_angle <= 19;
        242: s4_angle <= 20;
        243: s4_angle <= 22;
        244: s4_angle <= 23;
        245: s4_angle <= 24;
        246: s4_angle <= 26;
        247: s4_angle <= 27;
        248: s4_angle <= 28;
        249: s4_angle <= 29;
        250: s4_angle <= 30;
        251: s4_angle <= 31;
        252: s4_angle <= 0;
        253: s4_angle <= 2;
        254: s4_angle <= 4;
        255: s4_angle <= 5;
        256: s4_angle <= 7;
        257: s4_angle <= 9;
        258: s4_angle <= 10;
        259: s4_angle <= 12;
        260: s4_angle <= 14;
        261: s4_angle <= 15;
        262: s4_angle <= 17;
        263: s4_angle <= 18;
        264: s4_angle <= 20;
        265: s4_angle <= 21;
        266: s4_angle <= 22;
        267: s4_angle <= 24;
        268: s4_angle <= 25;
        269: s4_angle <= 26;
        270: s4_angle <= 27;
        271: s4_angle <= 28;
        272: s4_angle <= 29;
        273: s4_angle <= 30;
        274: s4_angle <= 31;
        275: s4_angle <= 0;
        276: s4_angle <= 2;
        277: s4_angle <= 3;
        278: s4_angle <= 5;
        279: s4_angle <= 7;
        280: s4_angle <= 8;
        281: s4_angle <= 10;
        282: s4_angle <= 12;
        283: s4_angle <= 13;
        284: s4_angle <= 15;
        285: s4_angle <= 16;
        286: s4_angle <= 18;
        287: s4_angle <= 19;
        288: s4_angle <= 20;
        289: s4_angle <= 22;
        290: s4_angle <= 23;
        291: s4_angle <= 24;
        292: s4_angle <= 25;
        293: s4_angle <= 26;
        294: s4_angle <= 27;
        295: s4_angle <= 28;
        296: s4_angle <= 29;
        297: s4_angle <= 30;
        298: s4_angle <= 31;
        299: s4_angle <= 0;
        300: s4_angle <= 2;
        301: s4_angle <= 3;
        302: s4_angle <= 5;
        303: s4_angle <= 6;
        304: s4_angle <= 8;
        305: s4_angle <= 10;
        306: s4_angle <= 11;
        307: s4_angle <= 13;
        308: s4_angle <= 14;
        309: s4_angle <= 16;
        310: s4_angle <= 17;
        311: s4_angle <= 18;
        312: s4_angle <= 20;
        313: s4_angle <= 21;
        314: s4_angle <= 22;
        315: s4_angle <= 23;
        316: s4_angle <= 24;
        317: s4_angle <= 25;
        318: s4_angle <= 26;
        319: s4_angle <= 27;
        320: s4_angle <= 28;
        321: s4_angle <= 29;
        322: s4_angle <= 30;
        323: s4_angle <= 31;
        324: s4_angle <= 0;
        325: s4_angle <= 2;
        326: s4_angle <= 3;
        327: s4_angle <= 5;
        328: s4_angle <= 6;
        329: s4_angle <= 8;
        330: s4_angle <= 9;
        331: s4_angle <= 11;
        332: s4_angle <= 12;
        333: s4_angle <= 14;
        334: s4_angle <= 15;
        335: s4_angle <= 16;
        336: s4_angle <= 18;
        337: s4_angle <= 19;
        338: s4_angle <= 20;
        339: s4_angle <= 21;
        340: s4_angle <= 22;
        341: s4_angle <= 24;
        342: s4_angle <= 25;
        343: s4_angle <= 26;
        344: s4_angle <= 27;
        345: s4_angle <= 28;
        346: s4_angle <= 29;
        347: s4_angle <= 30;
        348: s4_angle <= 30;
        349: s4_angle <= 31;
        350: s4_angle <= 0;
        351: s4_angle <= 2;
        352: s4_angle <= 3;
        353: s4_angle <= 5;
        354: s4_angle <= 6;
        355: s4_angle <= 7;
        356: s4_angle <= 9;
        357: s4_angle <= 10;
        358: s4_angle <= 12;
        359: s4_angle <= 13;
        360: s4_angle <= 14;
        361: s4_angle <= 16;
        362: s4_angle <= 17;
        363: s4_angle <= 18;
        364: s4_angle <= 19;
        365: s4_angle <= 21;
        366: s4_angle <= 22;
        367: s4_angle <= 23;
        368: s4_angle <= 24;
        369: s4_angle <= 25;
        370: s4_angle <= 26;
        371: s4_angle <= 27;
        372: s4_angle <= 28;
        373: s4_angle <= 29;
        374: s4_angle <= 30;
        375: s4_angle <= 30;
        376: s4_angle <= 31;
        377: s4_angle <= 0;
        378: s4_angle <= 1;
        379: s4_angle <= 3;
        380: s4_angle <= 4;
        381: s4_angle <= 6;
        382: s4_angle <= 7;
        383: s4_angle <= 9;
        384: s4_angle <= 10;
        385: s4_angle <= 11;
        386: s4_angle <= 13;
        387: s4_angle <= 14;
        388: s4_angle <= 15;
        389: s4_angle <= 16;
        390: s4_angle <= 18;
        391: s4_angle <= 19;
        392: s4_angle <= 20;
        393: s4_angle <= 21;
        394: s4_angle <= 22;
        395: s4_angle <= 23;
        396: s4_angle <= 24;
        397: s4_angle <= 25;
        398: s4_angle <= 26;
        399: s4_angle <= 27;
        400: s4_angle <= 28;
        401: s4_angle <= 29;
        402: s4_angle <= 30;
        403: s4_angle <= 30;
        404: s4_angle <= 31;
        405: s4_angle <= 0;
        406: s4_angle <= 1;
        407: s4_angle <= 3;
        408: s4_angle <= 4;
        409: s4_angle <= 6;
        410: s4_angle <= 7;
        411: s4_angle <= 8;
        412: s4_angle <= 10;
        413: s4_angle <= 11;
        414: s4_angle <= 12;
        415: s4_angle <= 14;
        416: s4_angle <= 15;
        417: s4_angle <= 16;
        418: s4_angle <= 17;
        419: s4_angle <= 18;
        420: s4_angle <= 19;
        421: s4_angle <= 21;
        422: s4_angle <= 22;
        423: s4_angle <= 23;
        424: s4_angle <= 24;
        425: s4_angle <= 25;
        426: s4_angle <= 26;
        427: s4_angle <= 26;
        428: s4_angle <= 27;
        429: s4_angle <= 28;
        430: s4_angle <= 29;
        431: s4_angle <= 30;
        432: s4_angle <= 31;
        433: s4_angle <= 31;
        434: s4_angle <= 0;
        435: s4_angle <= 1;
        436: s4_angle <= 3;
        437: s4_angle <= 4;
        438: s4_angle <= 5;
        439: s4_angle <= 7;
        440: s4_angle <= 8;
        441: s4_angle <= 9;
        442: s4_angle <= 11;
        443: s4_angle <= 12;
        444: s4_angle <= 13;
        445: s4_angle <= 14;
        446: s4_angle <= 16;
        447: s4_angle <= 17;
        448: s4_angle <= 18;
        449: s4_angle <= 19;
        450: s4_angle <= 20;
        451: s4_angle <= 21;
        452: s4_angle <= 22;
        453: s4_angle <= 23;
        454: s4_angle <= 24;
        455: s4_angle <= 25;
        456: s4_angle <= 26;
        457: s4_angle <= 27;
        458: s4_angle <= 27;
        459: s4_angle <= 28;
        460: s4_angle <= 29;
        461: s4_angle <= 30;
        462: s4_angle <= 31;
        463: s4_angle <= 31;
        464: s4_angle <= 0;
        465: s4_angle <= 1;
        466: s4_angle <= 3;
        467: s4_angle <= 4;
        468: s4_angle <= 5;
        469: s4_angle <= 7;
        470: s4_angle <= 8;
        471: s4_angle <= 9;
        472: s4_angle <= 10;
        473: s4_angle <= 12;
        474: s4_angle <= 13;
        475: s4_angle <= 14;
        476: s4_angle <= 15;
        477: s4_angle <= 16;
        478: s4_angle <= 17;
        479: s4_angle <= 18;
        480: s4_angle <= 19;
        481: s4_angle <= 20;
        482: s4_angle <= 21;
        483: s4_angle <= 22;
        484: s4_angle <= 23;
        485: s4_angle <= 24;
        486: s4_angle <= 25;
        487: s4_angle <= 26;
        488: s4_angle <= 27;
        489: s4_angle <= 28;
        490: s4_angle <= 28;
        491: s4_angle <= 29;
        492: s4_angle <= 30;
        493: s4_angle <= 31;
        494: s4_angle <= 31;
        495: s4_angle <= 0;
        496: s4_angle <= 1;
        497: s4_angle <= 3;
        498: s4_angle <= 4;
        499: s4_angle <= 5;
        500: s4_angle <= 6;
        501: s4_angle <= 8;
        502: s4_angle <= 9;
        503: s4_angle <= 10;
        504: s4_angle <= 11;
        505: s4_angle <= 12;
        506: s4_angle <= 13;
        507: s4_angle <= 15;
        508: s4_angle <= 16;
        509: s4_angle <= 17;
        510: s4_angle <= 18;
        511: s4_angle <= 19;
        512: s4_angle <= 20;
        513: s4_angle <= 21;
        514: s4_angle <= 22;
        515: s4_angle <= 23;
        516: s4_angle <= 24;
        517: s4_angle <= 25;
        518: s4_angle <= 25;
        519: s4_angle <= 26;
        520: s4_angle <= 27;
        521: s4_angle <= 28;
        522: s4_angle <= 29;
        523: s4_angle <= 29;
        524: s4_angle <= 30;
        525: s4_angle <= 31;
        526: s4_angle <= 31;
        527: s4_angle <= 0;
        528: s4_angle <= 1;
        529: s4_angle <= 2;
        530: s4_angle <= 4;
        531: s4_angle <= 5;
        532: s4_angle <= 6;
        533: s4_angle <= 7;
        534: s4_angle <= 9;
        535: s4_angle <= 10;
        536: s4_angle <= 11;
        537: s4_angle <= 12;
        538: s4_angle <= 13;
        539: s4_angle <= 14;
        540: s4_angle <= 15;
        541: s4_angle <= 16;
        542: s4_angle <= 17;
        543: s4_angle <= 18;
        544: s4_angle <= 19;
        545: s4_angle <= 20;
        546: s4_angle <= 21;
        547: s4_angle <= 22;
        548: s4_angle <= 23;
        549: s4_angle <= 24;
        550: s4_angle <= 25;
        551: s4_angle <= 26;
        552: s4_angle <= 26;
        553: s4_angle <= 27;
        554: s4_angle <= 28;
        555: s4_angle <= 29;
        556: s4_angle <= 29;
        557: s4_angle <= 30;
        558: s4_angle <= 31;
        559: s4_angle <= 31;
        560: s4_angle <= 0;
        561: s4_angle <= 1;
        562: s4_angle <= 2;
        563: s4_angle <= 4;
        564: s4_angle <= 5;
        565: s4_angle <= 6;
        566: s4_angle <= 7;
        567: s4_angle <= 8;
        568: s4_angle <= 9;
        569: s4_angle <= 11;
        570: s4_angle <= 12;
        571: s4_angle <= 13;
        572: s4_angle <= 14;
        573: s4_angle <= 15;
        574: s4_angle <= 16;
        575: s4_angle <= 17;
        576: s4_angle <= 18;
        577: s4_angle <= 19;
        578: s4_angle <= 20;
        579: s4_angle <= 21;
        580: s4_angle <= 22;
        581: s4_angle <= 23;
        582: s4_angle <= 23;
        583: s4_angle <= 24;
        584: s4_angle <= 25;
        585: s4_angle <= 26;
        586: s4_angle <= 27;
        587: s4_angle <= 27;
        588: s4_angle <= 28;
        589: s4_angle <= 29;
        590: s4_angle <= 29;
        591: s4_angle <= 30;
        592: s4_angle <= 31;
        593: s4_angle <= 31;
        594: s4_angle <= 0;
        595: s4_angle <= 1;
        596: s4_angle <= 2;
        597: s4_angle <= 3;
        598: s4_angle <= 5;
        599: s4_angle <= 6;
        600: s4_angle <= 7;
        601: s4_angle <= 8;
        602: s4_angle <= 9;
        603: s4_angle <= 10;
        604: s4_angle <= 11;
        605: s4_angle <= 12;
        606: s4_angle <= 13;
        607: s4_angle <= 14;
        608: s4_angle <= 16;
        609: s4_angle <= 16;
        610: s4_angle <= 17;
        611: s4_angle <= 18;
        612: s4_angle <= 19;
        613: s4_angle <= 20;
        614: s4_angle <= 21;
        615: s4_angle <= 22;
        616: s4_angle <= 23;
        617: s4_angle <= 24;
        618: s4_angle <= 24;
        619: s4_angle <= 25;
        620: s4_angle <= 26;
        621: s4_angle <= 27;
        622: s4_angle <= 27;
        623: s4_angle <= 28;
        624: s4_angle <= 29;
        625: s4_angle <= 30;
        626: s4_angle <= 30;
        627: s4_angle <= 31;
        628: s4_angle <= 31;
        629: s4_angle <= 0;
        630: s4_angle <= 1;
        631: s4_angle <= 2;
        632: s4_angle <= 3;
        633: s4_angle <= 5;
        634: s4_angle <= 6;
        635: s4_angle <= 7;
        636: s4_angle <= 8;
        637: s4_angle <= 9;
        638: s4_angle <= 10;
        639: s4_angle <= 11;
        640: s4_angle <= 12;
        641: s4_angle <= 13;
        642: s4_angle <= 14;
        643: s4_angle <= 15;
        644: s4_angle <= 16;
        645: s4_angle <= 17;
        646: s4_angle <= 18;
        647: s4_angle <= 19;
        648: s4_angle <= 20;
        649: s4_angle <= 21;
        650: s4_angle <= 22;
        651: s4_angle <= 22;
        652: s4_angle <= 23;
        653: s4_angle <= 24;
        654: s4_angle <= 25;
        655: s4_angle <= 25;
        656: s4_angle <= 26;
        657: s4_angle <= 27;
        658: s4_angle <= 28;
        659: s4_angle <= 28;
        660: s4_angle <= 29;
        661: s4_angle <= 30;
        662: s4_angle <= 30;
        663: s4_angle <= 31;
        664: s4_angle <= 31;
        665: s4_angle <= 0;
        666: s4_angle <= 1;
        667: s4_angle <= 2;
        668: s4_angle <= 3;
        669: s4_angle <= 4;
        670: s4_angle <= 5;
        671: s4_angle <= 7;
        672: s4_angle <= 8;
        673: s4_angle <= 9;
        674: s4_angle <= 10;
        675: s4_angle <= 11;
        676: s4_angle <= 12;
        677: s4_angle <= 13;
        678: s4_angle <= 14;
        679: s4_angle <= 15;
        680: s4_angle <= 16;
        681: s4_angle <= 17;
        682: s4_angle <= 18;
        683: s4_angle <= 18;
        684: s4_angle <= 19;
        685: s4_angle <= 20;
        686: s4_angle <= 21;
        687: s4_angle <= 22;
        688: s4_angle <= 23;
        689: s4_angle <= 23;
        690: s4_angle <= 24;
        691: s4_angle <= 25;
        692: s4_angle <= 26;
        693: s4_angle <= 26;
        694: s4_angle <= 27;
        695: s4_angle <= 28;
        696: s4_angle <= 28;
        697: s4_angle <= 29;
        698: s4_angle <= 30;
        699: s4_angle <= 30;
        700: s4_angle <= 31;
        701: s4_angle <= 31;
        702: s4_angle <= 0;
        703: s4_angle <= 1;
        704: s4_angle <= 2;
        705: s4_angle <= 3;
        706: s4_angle <= 4;
        707: s4_angle <= 5;
        708: s4_angle <= 6;
        709: s4_angle <= 7;
        710: s4_angle <= 8;
        711: s4_angle <= 9;
        712: s4_angle <= 10;
        713: s4_angle <= 11;
        714: s4_angle <= 12;
        715: s4_angle <= 13;
        716: s4_angle <= 14;
        717: s4_angle <= 15;
        718: s4_angle <= 16;
        719: s4_angle <= 17;
        720: s4_angle <= 18;
        721: s4_angle <= 19;
        722: s4_angle <= 20;
        723: s4_angle <= 21;
        724: s4_angle <= 21;
        725: s4_angle <= 22;
        726: s4_angle <= 23;
        727: s4_angle <= 24;
        728: s4_angle <= 24;
        729: s4_angle <= 25;
        730: s4_angle <= 26;
        731: s4_angle <= 27;
        732: s4_angle <= 27;
        733: s4_angle <= 28;
        734: s4_angle <= 29;
        735: s4_angle <= 29;
        736: s4_angle <= 30;
        737: s4_angle <= 30;
        738: s4_angle <= 31;
        739: s4_angle <= 31;
        740: s4_angle <= 0;
        741: s4_angle <= 1;
        742: s4_angle <= 2;
        743: s4_angle <= 3;
        744: s4_angle <= 4;
        745: s4_angle <= 5;
        746: s4_angle <= 6;
        747: s4_angle <= 7;
        748: s4_angle <= 8;
        749: s4_angle <= 9;
        750: s4_angle <= 10;
        751: s4_angle <= 11;
        752: s4_angle <= 12;
        753: s4_angle <= 13;
        754: s4_angle <= 14;
        755: s4_angle <= 15;
        756: s4_angle <= 16;
        757: s4_angle <= 17;
        758: s4_angle <= 18;
        759: s4_angle <= 18;
        760: s4_angle <= 19;
        761: s4_angle <= 20;
        762: s4_angle <= 21;
        763: s4_angle <= 22;
        764: s4_angle <= 22;
        765: s4_angle <= 23;
        766: s4_angle <= 24;
        767: s4_angle <= 25;
        768: s4_angle <= 25;
        769: s4_angle <= 26;
        770: s4_angle <= 27;
        771: s4_angle <= 27;
        772: s4_angle <= 28;
        773: s4_angle <= 29;
        774: s4_angle <= 29;
        775: s4_angle <= 30;
        776: s4_angle <= 30;
        777: s4_angle <= 31;
        778: s4_angle <= 31;
        779: s4_angle <= 0;
        780: s4_angle <= 1;
        781: s4_angle <= 2;
        782: s4_angle <= 3;
        783: s4_angle <= 4;
        784: s4_angle <= 5;
        785: s4_angle <= 6;
        786: s4_angle <= 7;
        787: s4_angle <= 8;
        788: s4_angle <= 9;
        789: s4_angle <= 10;
        790: s4_angle <= 11;
        791: s4_angle <= 12;
        792: s4_angle <= 13;
        793: s4_angle <= 14;
        794: s4_angle <= 15;
        795: s4_angle <= 16;
        796: s4_angle <= 16;
        797: s4_angle <= 17;
        798: s4_angle <= 18;
        799: s4_angle <= 19;
        800: s4_angle <= 20;
        801: s4_angle <= 20;
        802: s4_angle <= 21;
        803: s4_angle <= 22;
        804: s4_angle <= 23;
        805: s4_angle <= 23;
        806: s4_angle <= 24;
        807: s4_angle <= 25;
        808: s4_angle <= 26;
        809: s4_angle <= 26;
        810: s4_angle <= 27;
        811: s4_angle <= 27;
        812: s4_angle <= 28;
        813: s4_angle <= 29;
        814: s4_angle <= 29;
        815: s4_angle <= 30;
        816: s4_angle <= 30;
        817: s4_angle <= 31;
        818: s4_angle <= 31;
        819: s4_angle <= 0;
        820: s4_angle <= 1;
        821: s4_angle <= 2;
        822: s4_angle <= 3;
        823: s4_angle <= 4;
        824: s4_angle <= 5;
        825: s4_angle <= 6;
        826: s4_angle <= 7;
        827: s4_angle <= 8;
        828: s4_angle <= 9;
        829: s4_angle <= 10;
        830: s4_angle <= 11;
        831: s4_angle <= 12;
        832: s4_angle <= 13;
        833: s4_angle <= 13;
        834: s4_angle <= 14;
        835: s4_angle <= 15;
        836: s4_angle <= 16;
        837: s4_angle <= 17;
        838: s4_angle <= 18;
        839: s4_angle <= 18;
        840: s4_angle <= 19;
        841: s4_angle <= 20;
        842: s4_angle <= 21;
        843: s4_angle <= 22;
        844: s4_angle <= 22;
        845: s4_angle <= 23;
        846: s4_angle <= 24;
        847: s4_angle <= 24;
        848: s4_angle <= 25;
        849: s4_angle <= 26;
        850: s4_angle <= 26;
        851: s4_angle <= 27;
        852: s4_angle <= 28;
        853: s4_angle <= 28;
        854: s4_angle <= 29;
        855: s4_angle <= 29;
        856: s4_angle <= 30;
        857: s4_angle <= 30;
        858: s4_angle <= 31;
        859: s4_angle <= 31;
        860: s4_angle <= 0;
        861: s4_angle <= 1;
        862: s4_angle <= 2;
        863: s4_angle <= 3;
        864: s4_angle <= 4;
        865: s4_angle <= 5;
        866: s4_angle <= 6;
        867: s4_angle <= 7;
        868: s4_angle <= 8;
        869: s4_angle <= 9;
        870: s4_angle <= 10;
        871: s4_angle <= 10;
        872: s4_angle <= 11;
        873: s4_angle <= 12;
        874: s4_angle <= 13;
        875: s4_angle <= 14;
        876: s4_angle <= 15;
        877: s4_angle <= 16;
        878: s4_angle <= 16;
        879: s4_angle <= 17;
        880: s4_angle <= 18;
        881: s4_angle <= 19;
        882: s4_angle <= 20;
        883: s4_angle <= 20;
        884: s4_angle <= 21;
        885: s4_angle <= 22;
        886: s4_angle <= 23;
        887: s4_angle <= 23;
        888: s4_angle <= 24;
        889: s4_angle <= 25;
        890: s4_angle <= 25;
        891: s4_angle <= 26;
        892: s4_angle <= 27;
        893: s4_angle <= 27;
        894: s4_angle <= 28;
        895: s4_angle <= 28;
        896: s4_angle <= 29;
        897: s4_angle <= 29;
        898: s4_angle <= 30;
        899: s4_angle <= 30;
        900: s4_angle <= 31;
        901: s4_angle <= 31;
        902: s4_angle <= 0;
        903: s4_angle <= 1;
        904: s4_angle <= 2;
        905: s4_angle <= 3;
        906: s4_angle <= 4;
        907: s4_angle <= 5;
        908: s4_angle <= 6;
        909: s4_angle <= 7;
        910: s4_angle <= 7;
        911: s4_angle <= 8;
        912: s4_angle <= 9;
        913: s4_angle <= 10;
        914: s4_angle <= 11;
        915: s4_angle <= 12;
        916: s4_angle <= 13;
        917: s4_angle <= 14;
        918: s4_angle <= 15;
        919: s4_angle <= 15;
        920: s4_angle <= 16;
        921: s4_angle <= 17;
        922: s4_angle <= 18;
        923: s4_angle <= 19;
        924: s4_angle <= 19;
        925: s4_angle <= 20;
        926: s4_angle <= 21;
        927: s4_angle <= 21;
        928: s4_angle <= 22;
        929: s4_angle <= 23;
        930: s4_angle <= 24;
        931: s4_angle <= 24;
        932: s4_angle <= 25;
        933: s4_angle <= 25;
        934: s4_angle <= 26;
        935: s4_angle <= 27;
        936: s4_angle <= 27;
        937: s4_angle <= 28;
        938: s4_angle <= 28;
        939: s4_angle <= 29;
        940: s4_angle <= 29;
        941: s4_angle <= 30;
        942: s4_angle <= 31;
        943: s4_angle <= 31;
        944: s4_angle <= 31;
        945: s4_angle <= 0;
        946: s4_angle <= 1;
        947: s4_angle <= 2;
        948: s4_angle <= 3;
        949: s4_angle <= 4;
        950: s4_angle <= 5;
        951: s4_angle <= 6;
        952: s4_angle <= 6;
        953: s4_angle <= 7;
        954: s4_angle <= 8;
        955: s4_angle <= 9;
        956: s4_angle <= 10;
        957: s4_angle <= 11;
        958: s4_angle <= 12;
        959: s4_angle <= 13;
        960: s4_angle <= 13;
        961: s4_angle <= 14;
        962: s4_angle <= 15;
        963: s4_angle <= 16;
        964: s4_angle <= 17;
        965: s4_angle <= 17;
        966: s4_angle <= 18;
        967: s4_angle <= 19;
        968: s4_angle <= 20;
        969: s4_angle <= 20;
        970: s4_angle <= 21;
        971: s4_angle <= 22;
        972: s4_angle <= 22;
        973: s4_angle <= 23;
        974: s4_angle <= 24;
        975: s4_angle <= 24;
        976: s4_angle <= 25;
        977: s4_angle <= 26;
        978: s4_angle <= 26;
        979: s4_angle <= 27;
        980: s4_angle <= 27;
        981: s4_angle <= 28;
        982: s4_angle <= 28;
        983: s4_angle <= 29;
        984: s4_angle <= 30;
        985: s4_angle <= 30;
        986: s4_angle <= 31;
        987: s4_angle <= 31;
        988: s4_angle <= 31;
        989: s4_angle <= 0;
        990: s4_angle <= 1;
        991: s4_angle <= 2;
        992: s4_angle <= 3;
        993: s4_angle <= 4;
        994: s4_angle <= 5;
        995: s4_angle <= 5;
        996: s4_angle <= 6;
        997: s4_angle <= 7;
        998: s4_angle <= 8;
        999: s4_angle <= 9;
        1000: s4_angle <= 10;
        1001: s4_angle <= 11;
        1002: s4_angle <= 11;
        1003: s4_angle <= 12;
        1004: s4_angle <= 13;
        1005: s4_angle <= 14;
        1006: s4_angle <= 15;
        1007: s4_angle <= 16;
        1008: s4_angle <= 16;
        1009: s4_angle <= 17;
        1010: s4_angle <= 18;
        1011: s4_angle <= 19;
        1012: s4_angle <= 19;
        1013: s4_angle <= 20;
        1014: s4_angle <= 21;
        1015: s4_angle <= 21;
        1016: s4_angle <= 22;
        1017: s4_angle <= 23;
        1018: s4_angle <= 23;
        1019: s4_angle <= 24;
        1020: s4_angle <= 25;
        1021: s4_angle <= 25;
        1022: s4_angle <= 26;
        1023: s4_angle <= 26;
        1024: s4_angle <= 27;
        1025: s4_angle <= 27;
        1026: s4_angle <= 28;
        1027: s4_angle <= 29;
        1028: s4_angle <= 29;
        1029: s4_angle <= 30;
        1030: s4_angle <= 30;
        1031: s4_angle <= 31;
        1032: s4_angle <= 31;
        1033: s4_angle <= 31;
        1034: s4_angle <= 0;
        1035: s4_angle <= 1;
        1036: s4_angle <= 2;
        1037: s4_angle <= 3;
        1038: s4_angle <= 4;
        1039: s4_angle <= 4;
        1040: s4_angle <= 5;
        1041: s4_angle <= 6;
        1042: s4_angle <= 7;
        1043: s4_angle <= 8;
        1044: s4_angle <= 9;
        1045: s4_angle <= 10;
        1046: s4_angle <= 10;
        1047: s4_angle <= 11;
        1048: s4_angle <= 12;
        1049: s4_angle <= 13;
        1050: s4_angle <= 14;
        1051: s4_angle <= 14;
        1052: s4_angle <= 15;
        1053: s4_angle <= 16;
        1054: s4_angle <= 17;
        1055: s4_angle <= 17;
        1056: s4_angle <= 18;
        1057: s4_angle <= 19;
        1058: s4_angle <= 20;
        1059: s4_angle <= 20;
        1060: s4_angle <= 21;
        1061: s4_angle <= 22;
        1062: s4_angle <= 22;
        1063: s4_angle <= 23;
        1064: s4_angle <= 24;
        1065: s4_angle <= 24;
        1066: s4_angle <= 25;
        1067: s4_angle <= 25;
        1068: s4_angle <= 26;
        1069: s4_angle <= 27;
        1070: s4_angle <= 27;
        1071: s4_angle <= 28;
        1072: s4_angle <= 28;
        1073: s4_angle <= 29;
        1074: s4_angle <= 29;
        1075: s4_angle <= 30;
        1076: s4_angle <= 30;
        1077: s4_angle <= 31;
        1078: s4_angle <= 31;
        1079: s4_angle <= 31;
        1080: s4_angle <= 0;
        1081: s4_angle <= 1;
        1082: s4_angle <= 2;
        1083: s4_angle <= 3;
        1084: s4_angle <= 3;
        1085: s4_angle <= 4;
        1086: s4_angle <= 5;
        1087: s4_angle <= 6;
        1088: s4_angle <= 7;
        1089: s4_angle <= 8;
        1090: s4_angle <= 9;
        1091: s4_angle <= 9;
        1092: s4_angle <= 10;
        1093: s4_angle <= 11;
        1094: s4_angle <= 12;
        1095: s4_angle <= 13;
        1096: s4_angle <= 13;
        1097: s4_angle <= 14;
        1098: s4_angle <= 15;
        1099: s4_angle <= 16;
        1100: s4_angle <= 16;
        1101: s4_angle <= 17;
        1102: s4_angle <= 18;
        1103: s4_angle <= 19;
        1104: s4_angle <= 19;
        1105: s4_angle <= 20;
        1106: s4_angle <= 21;
        1107: s4_angle <= 21;
        1108: s4_angle <= 22;
        1109: s4_angle <= 23;
        1110: s4_angle <= 23;
        1111: s4_angle <= 24;
        1112: s4_angle <= 24;
        1113: s4_angle <= 25;
        1114: s4_angle <= 26;
        1115: s4_angle <= 26;
        1116: s4_angle <= 27;
        1117: s4_angle <= 27;
        1118: s4_angle <= 28;
        1119: s4_angle <= 28;
        1120: s4_angle <= 29;
        1121: s4_angle <= 29;
        1122: s4_angle <= 30;
        1123: s4_angle <= 30;
        1124: s4_angle <= 31;
        1125: s4_angle <= 31;
        1126: s4_angle <= 31;
        1127: s4_angle <= 0;
        1128: s4_angle <= 1;
        1129: s4_angle <= 2;
        1130: s4_angle <= 3;
        1131: s4_angle <= 3;
        1132: s4_angle <= 4;
        1133: s4_angle <= 5;
        1134: s4_angle <= 6;
        1135: s4_angle <= 7;
        1136: s4_angle <= 8;
        1137: s4_angle <= 8;
        1138: s4_angle <= 9;
        1139: s4_angle <= 10;
        1140: s4_angle <= 11;
        1141: s4_angle <= 12;
        1142: s4_angle <= 12;
        1143: s4_angle <= 13;
        1144: s4_angle <= 14;
        1145: s4_angle <= 15;
        1146: s4_angle <= 15;
        1147: s4_angle <= 16;
        1148: s4_angle <= 17;
        1149: s4_angle <= 18;
        1150: s4_angle <= 18;
        1151: s4_angle <= 19;
        1152: s4_angle <= 20;
        1153: s4_angle <= 20;
        1154: s4_angle <= 21;
        1155: s4_angle <= 22;
        1156: s4_angle <= 22;
        1157: s4_angle <= 23;
        1158: s4_angle <= 23;
        1159: s4_angle <= 24;
        1160: s4_angle <= 25;
        1161: s4_angle <= 25;
        1162: s4_angle <= 26;
        1163: s4_angle <= 26;
        1164: s4_angle <= 27;
        1165: s4_angle <= 27;
        1166: s4_angle <= 28;
        1167: s4_angle <= 28;
        1168: s4_angle <= 29;
        1169: s4_angle <= 29;
        1170: s4_angle <= 30;
        1171: s4_angle <= 30;
        1172: s4_angle <= 31;
        1173: s4_angle <= 31;
        1174: s4_angle <= 31;
        1175: s4_angle <= 0;
        1176: s4_angle <= 1;
        1177: s4_angle <= 2;
        1178: s4_angle <= 2;
        1179: s4_angle <= 3;
        1180: s4_angle <= 4;
        1181: s4_angle <= 5;
        1182: s4_angle <= 6;
        1183: s4_angle <= 7;
        1184: s4_angle <= 7;
        1185: s4_angle <= 8;
        1186: s4_angle <= 9;
        1187: s4_angle <= 10;
        1188: s4_angle <= 11;
        1189: s4_angle <= 11;
        1190: s4_angle <= 12;
        1191: s4_angle <= 13;
        1192: s4_angle <= 14;
        1193: s4_angle <= 14;
        1194: s4_angle <= 15;
        1195: s4_angle <= 16;
        1196: s4_angle <= 16;
        1197: s4_angle <= 17;
        1198: s4_angle <= 18;
        1199: s4_angle <= 19;
        1200: s4_angle <= 19;
        1201: s4_angle <= 20;
        1202: s4_angle <= 21;
        1203: s4_angle <= 21;
        1204: s4_angle <= 22;
        1205: s4_angle <= 22;
        1206: s4_angle <= 23;
        1207: s4_angle <= 24;
        1208: s4_angle <= 24;
        1209: s4_angle <= 25;
        1210: s4_angle <= 25;
        1211: s4_angle <= 26;
        1212: s4_angle <= 26;
        1213: s4_angle <= 27;
        1214: s4_angle <= 27;
        1215: s4_angle <= 28;
        1216: s4_angle <= 28;
        1217: s4_angle <= 29;
        1218: s4_angle <= 29;
        1219: s4_angle <= 30;
        1220: s4_angle <= 30;
        1221: s4_angle <= 31;
        1222: s4_angle <= 31;
        1223: s4_angle <= 31;
        1224: s4_angle <= 0;
        1225: s4_angle <= 1;
        1226: s4_angle <= 2;
        1227: s4_angle <= 2;
        1228: s4_angle <= 3;
        1229: s4_angle <= 4;
        1230: s4_angle <= 5;
        1231: s4_angle <= 6;
        1232: s4_angle <= 6;
        1233: s4_angle <= 7;
        1234: s4_angle <= 8;
        1235: s4_angle <= 9;
        1236: s4_angle <= 10;
        1237: s4_angle <= 10;
        1238: s4_angle <= 11;
        1239: s4_angle <= 12;
        1240: s4_angle <= 13;
        1241: s4_angle <= 13;
        1242: s4_angle <= 14;
        1243: s4_angle <= 15;
        1244: s4_angle <= 16;
        1245: s4_angle <= 16;
        1246: s4_angle <= 17;
        1247: s4_angle <= 18;
        1248: s4_angle <= 18;
        1249: s4_angle <= 19;
        1250: s4_angle <= 20;
        1251: s4_angle <= 20;
        1252: s4_angle <= 21;
        1253: s4_angle <= 21;
        1254: s4_angle <= 22;
        1255: s4_angle <= 23;
        1256: s4_angle <= 23;
        1257: s4_angle <= 24;
        1258: s4_angle <= 24;
        1259: s4_angle <= 25;
        1260: s4_angle <= 25;
        1261: s4_angle <= 26;
        1262: s4_angle <= 26;
        1263: s4_angle <= 27;
        1264: s4_angle <= 27;
        1265: s4_angle <= 28;
        1266: s4_angle <= 28;
        1267: s4_angle <= 29;
        1268: s4_angle <= 29;
        1269: s4_angle <= 30;
        1270: s4_angle <= 30;
        1271: s4_angle <= 31;
        1272: s4_angle <= 31;
        1273: s4_angle <= 31;
        1274: s4_angle <= 0;
        1275: s4_angle <= 1;
        1276: s4_angle <= 2;
        1277: s4_angle <= 2;
        1278: s4_angle <= 3;
        1279: s4_angle <= 4;
        1280: s4_angle <= 5;
        1281: s4_angle <= 6;
        1282: s4_angle <= 6;
        1283: s4_angle <= 7;
        1284: s4_angle <= 8;
        1285: s4_angle <= 9;
        1286: s4_angle <= 9;
        1287: s4_angle <= 10;
        1288: s4_angle <= 11;
        1289: s4_angle <= 12;
        1290: s4_angle <= 12;
        1291: s4_angle <= 13;
        1292: s4_angle <= 14;
        1293: s4_angle <= 15;
        1294: s4_angle <= 15;
        1295: s4_angle <= 16;
        1296: s4_angle <= 17;
        1297: s4_angle <= 17;
        1298: s4_angle <= 18;
        1299: s4_angle <= 19;
        1300: s4_angle <= 19;
        1301: s4_angle <= 20;
        1302: s4_angle <= 20;
        1303: s4_angle <= 21;
        1304: s4_angle <= 22;
        1305: s4_angle <= 22;
        1306: s4_angle <= 23;
        1307: s4_angle <= 23;
        1308: s4_angle <= 24;
        1309: s4_angle <= 25;
        1310: s4_angle <= 25;
        1311: s4_angle <= 26;
        1312: s4_angle <= 26;
        1313: s4_angle <= 27;
        1314: s4_angle <= 27;
        1315: s4_angle <= 28;
        1316: s4_angle <= 28;
        1317: s4_angle <= 29;
        1318: s4_angle <= 29;
        1319: s4_angle <= 29;
        1320: s4_angle <= 30;
        1321: s4_angle <= 30;
        1322: s4_angle <= 31;
        1323: s4_angle <= 31;
        1324: s4_angle <= 31;
        1325: s4_angle <= 0;
        1326: s4_angle <= 1;
        1327: s4_angle <= 2;
        1328: s4_angle <= 2;
        1329: s4_angle <= 3;
        1330: s4_angle <= 4;
        1331: s4_angle <= 5;
        1332: s4_angle <= 5;
        1333: s4_angle <= 6;
        1334: s4_angle <= 7;
        1335: s4_angle <= 8;
        1336: s4_angle <= 8;
        1337: s4_angle <= 9;
        1338: s4_angle <= 10;
        1339: s4_angle <= 11;
        1340: s4_angle <= 11;
        1341: s4_angle <= 12;
        1342: s4_angle <= 13;
        1343: s4_angle <= 14;
        1344: s4_angle <= 14;
        1345: s4_angle <= 15;
        1346: s4_angle <= 16;
        1347: s4_angle <= 16;
        1348: s4_angle <= 17;
        1349: s4_angle <= 18;
        1350: s4_angle <= 18;
        1351: s4_angle <= 19;
        1352: s4_angle <= 20;
        1353: s4_angle <= 20;
        1354: s4_angle <= 21;
        1355: s4_angle <= 21;
        1356: s4_angle <= 22;
        1357: s4_angle <= 22;
        1358: s4_angle <= 23;
        1359: s4_angle <= 24;
        1360: s4_angle <= 24;
        1361: s4_angle <= 25;
        1362: s4_angle <= 25;
        1363: s4_angle <= 26;
        1364: s4_angle <= 26;
        1365: s4_angle <= 27;
        1366: s4_angle <= 27;
        1367: s4_angle <= 28;
        1368: s4_angle <= 28;
        1369: s4_angle <= 29;
        1370: s4_angle <= 29;
        1371: s4_angle <= 30;
        1372: s4_angle <= 30;
        1373: s4_angle <= 30;
        1374: s4_angle <= 31;
        1375: s4_angle <= 31;
        1376: s4_angle <= 31;
        1377: s4_angle <= 0;
        1378: s4_angle <= 1;
        1379: s4_angle <= 2;
        1380: s4_angle <= 2;
        1381: s4_angle <= 3;
        1382: s4_angle <= 4;
        1383: s4_angle <= 5;
        1384: s4_angle <= 5;
        1385: s4_angle <= 6;
        1386: s4_angle <= 7;
        1387: s4_angle <= 8;
        1388: s4_angle <= 8;
        1389: s4_angle <= 9;
        1390: s4_angle <= 10;
        1391: s4_angle <= 11;
        1392: s4_angle <= 11;
        1393: s4_angle <= 12;
        1394: s4_angle <= 13;
        1395: s4_angle <= 13;
        1396: s4_angle <= 14;
        1397: s4_angle <= 15;
        1398: s4_angle <= 15;
        1399: s4_angle <= 16;
        1400: s4_angle <= 17;
        1401: s4_angle <= 17;
        1402: s4_angle <= 18;
        1403: s4_angle <= 19;
        1404: s4_angle <= 19;
        1405: s4_angle <= 20;
        1406: s4_angle <= 20;
        1407: s4_angle <= 21;
        1408: s4_angle <= 22;
        1409: s4_angle <= 22;
        1410: s4_angle <= 23;
        1411: s4_angle <= 23;
        1412: s4_angle <= 24;
        1413: s4_angle <= 24;
        1414: s4_angle <= 25;
        1415: s4_angle <= 25;
        1416: s4_angle <= 26;
        1417: s4_angle <= 26;
        1418: s4_angle <= 27;
        1419: s4_angle <= 27;
        1420: s4_angle <= 28;
        1421: s4_angle <= 28;
        1422: s4_angle <= 29;
        1423: s4_angle <= 29;
        1424: s4_angle <= 30;
        1425: s4_angle <= 30;
        1426: s4_angle <= 30;
        1427: s4_angle <= 31;
        1428: s4_angle <= 31;
        1429: s4_angle <= 31;
        1430: s4_angle <= 0;
        1431: s4_angle <= 1;
        1432: s4_angle <= 2;
        1433: s4_angle <= 2;
        1434: s4_angle <= 3;
        1435: s4_angle <= 4;
        1436: s4_angle <= 5;
        1437: s4_angle <= 5;
        1438: s4_angle <= 6;
        1439: s4_angle <= 7;
        1440: s4_angle <= 7;
        1441: s4_angle <= 8;
        1442: s4_angle <= 9;
        1443: s4_angle <= 10;
        1444: s4_angle <= 10;
        1445: s4_angle <= 11;
        1446: s4_angle <= 12;
        1447: s4_angle <= 12;
        1448: s4_angle <= 13;
        1449: s4_angle <= 14;
        1450: s4_angle <= 14;
        1451: s4_angle <= 15;
        1452: s4_angle <= 16;
        1453: s4_angle <= 16;
        1454: s4_angle <= 17;
        1455: s4_angle <= 18;
        1456: s4_angle <= 18;
        1457: s4_angle <= 19;
        1458: s4_angle <= 19;
        1459: s4_angle <= 20;
        1460: s4_angle <= 21;
        1461: s4_angle <= 21;
        1462: s4_angle <= 22;
        1463: s4_angle <= 22;
        1464: s4_angle <= 23;
        1465: s4_angle <= 23;
        1466: s4_angle <= 24;
        1467: s4_angle <= 24;
        1468: s4_angle <= 25;
        1469: s4_angle <= 25;
        1470: s4_angle <= 26;
        1471: s4_angle <= 26;
        1472: s4_angle <= 27;
        1473: s4_angle <= 27;
        1474: s4_angle <= 28;
        1475: s4_angle <= 28;
        1476: s4_angle <= 29;
        1477: s4_angle <= 29;
        1478: s4_angle <= 30;
        1479: s4_angle <= 30;
        1480: s4_angle <= 30;
        1481: s4_angle <= 31;
        1482: s4_angle <= 31;
        1483: s4_angle <= 31;
        1484: s4_angle <= 0;
        1485: s4_angle <= 1;
        1486: s4_angle <= 1;
        1487: s4_angle <= 2;
        1488: s4_angle <= 3;
        1489: s4_angle <= 4;
        1490: s4_angle <= 4;
        1491: s4_angle <= 5;
        1492: s4_angle <= 6;
        1493: s4_angle <= 7;
        1494: s4_angle <= 7;
        1495: s4_angle <= 8;
        1496: s4_angle <= 9;
        1497: s4_angle <= 9;
        1498: s4_angle <= 10;
        1499: s4_angle <= 11;
        1500: s4_angle <= 12;
        1501: s4_angle <= 12;
        1502: s4_angle <= 13;
        1503: s4_angle <= 14;
        1504: s4_angle <= 14;
        1505: s4_angle <= 15;
        1506: s4_angle <= 16;
        1507: s4_angle <= 16;
        1508: s4_angle <= 17;
        1509: s4_angle <= 17;
        1510: s4_angle <= 18;
        1511: s4_angle <= 19;
        1512: s4_angle <= 19;
        1513: s4_angle <= 20;
        1514: s4_angle <= 20;
        1515: s4_angle <= 21;
        1516: s4_angle <= 21;
        1517: s4_angle <= 22;
        1518: s4_angle <= 23;
        1519: s4_angle <= 23;
        1520: s4_angle <= 24;
        1521: s4_angle <= 24;
        1522: s4_angle <= 25;
        1523: s4_angle <= 25;
        1524: s4_angle <= 26;
        1525: s4_angle <= 26;
        1526: s4_angle <= 27;
        1527: s4_angle <= 27;
        1528: s4_angle <= 27;
        1529: s4_angle <= 28;
        1530: s4_angle <= 28;
        1531: s4_angle <= 29;
        1532: s4_angle <= 29;
        1533: s4_angle <= 30;
        1534: s4_angle <= 30;
        1535: s4_angle <= 30;
        1536: s4_angle <= 31;
        1537: s4_angle <= 31;
        1538: s4_angle <= 31;
        1539: s4_angle <= 0;
        1540: s4_angle <= 1;
        1541: s4_angle <= 1;
        1542: s4_angle <= 2;
        1543: s4_angle <= 3;
        1544: s4_angle <= 4;
        1545: s4_angle <= 4;
        1546: s4_angle <= 5;
        1547: s4_angle <= 6;
        1548: s4_angle <= 6;
        1549: s4_angle <= 7;
        1550: s4_angle <= 8;
        1551: s4_angle <= 9;
        1552: s4_angle <= 9;
        1553: s4_angle <= 10;
        1554: s4_angle <= 11;
        1555: s4_angle <= 11;
        1556: s4_angle <= 12;
        1557: s4_angle <= 13;
        1558: s4_angle <= 13;
        1559: s4_angle <= 14;
        1560: s4_angle <= 15;
        1561: s4_angle <= 15;
        1562: s4_angle <= 16;
        1563: s4_angle <= 16;
        1564: s4_angle <= 17;
        1565: s4_angle <= 18;
        1566: s4_angle <= 18;
        1567: s4_angle <= 19;
        1568: s4_angle <= 19;
        1569: s4_angle <= 20;
        1570: s4_angle <= 21;
        1571: s4_angle <= 21;
        1572: s4_angle <= 22;
        1573: s4_angle <= 22;
        1574: s4_angle <= 23;
        1575: s4_angle <= 23;
        1576: s4_angle <= 24;
        1577: s4_angle <= 24;
        1578: s4_angle <= 25;
        1579: s4_angle <= 25;
        1580: s4_angle <= 26;
        1581: s4_angle <= 26;
        1582: s4_angle <= 27;
        1583: s4_angle <= 27;
        1584: s4_angle <= 28;
        1585: s4_angle <= 28;
        1586: s4_angle <= 28;
        1587: s4_angle <= 29;
        1588: s4_angle <= 29;
        1589: s4_angle <= 30;
        1590: s4_angle <= 30;
        1591: s4_angle <= 30;
        1592: s4_angle <= 31;
        1593: s4_angle <= 31;
        1594: s4_angle <= 31;
        1595: s4_angle <= 0;
        1596: s4_angle <= 1;
        1597: s4_angle <= 1;
        1598: s4_angle <= 2;
        1599: s4_angle <= 3;
        1600: s4_angle <= 4;
        1601: s4_angle <= 4;
        1602: s4_angle <= 5;
        1603: s4_angle <= 6;
        1604: s4_angle <= 6;
        1605: s4_angle <= 7;
        1606: s4_angle <= 8;
        1607: s4_angle <= 8;
        1608: s4_angle <= 9;
        1609: s4_angle <= 10;
        1610: s4_angle <= 10;
        1611: s4_angle <= 11;
        1612: s4_angle <= 12;
        1613: s4_angle <= 12;
        1614: s4_angle <= 13;
        1615: s4_angle <= 14;
        1616: s4_angle <= 14;
        1617: s4_angle <= 15;
        1618: s4_angle <= 16;
        1619: s4_angle <= 16;
        1620: s4_angle <= 17;
        1621: s4_angle <= 17;
        1622: s4_angle <= 18;
        1623: s4_angle <= 19;
        1624: s4_angle <= 19;
        1625: s4_angle <= 20;
        1626: s4_angle <= 20;
        1627: s4_angle <= 21;
        1628: s4_angle <= 21;
        1629: s4_angle <= 22;
        1630: s4_angle <= 22;
        1631: s4_angle <= 23;
        1632: s4_angle <= 23;
        1633: s4_angle <= 24;
        1634: s4_angle <= 24;
        1635: s4_angle <= 25;
        1636: s4_angle <= 25;
        1637: s4_angle <= 26;
        1638: s4_angle <= 26;
        1639: s4_angle <= 27;
        1640: s4_angle <= 27;
        1641: s4_angle <= 28;
        1642: s4_angle <= 28;
        1643: s4_angle <= 29;
        1644: s4_angle <= 29;
        1645: s4_angle <= 29;
        1646: s4_angle <= 30;
        1647: s4_angle <= 30;
        1648: s4_angle <= 31;
        1649: s4_angle <= 31;
        1650: s4_angle <= 31;
        1651: s4_angle <= 31;
        1652: s4_angle <= 0;
        1653: s4_angle <= 1;
        1654: s4_angle <= 1;
        1655: s4_angle <= 2;
        1656: s4_angle <= 3;
        1657: s4_angle <= 4;
        1658: s4_angle <= 4;
        1659: s4_angle <= 5;
        1660: s4_angle <= 6;
        1661: s4_angle <= 6;
        1662: s4_angle <= 7;
        1663: s4_angle <= 8;
        1664: s4_angle <= 8;
        1665: s4_angle <= 9;
        1666: s4_angle <= 10;
        1667: s4_angle <= 10;
        1668: s4_angle <= 11;
        1669: s4_angle <= 12;
        1670: s4_angle <= 12;
        1671: s4_angle <= 13;
        1672: s4_angle <= 14;
        1673: s4_angle <= 14;
        1674: s4_angle <= 15;
        1675: s4_angle <= 15;
        1676: s4_angle <= 16;
        1677: s4_angle <= 17;
        1678: s4_angle <= 17;
        1679: s4_angle <= 18;
        1680: s4_angle <= 18;
        1681: s4_angle <= 19;
        1682: s4_angle <= 19;
        1683: s4_angle <= 20;
        1684: s4_angle <= 21;
        1685: s4_angle <= 21;
        1686: s4_angle <= 22;
        1687: s4_angle <= 22;
        1688: s4_angle <= 23;
        1689: s4_angle <= 23;
        1690: s4_angle <= 24;
        1691: s4_angle <= 24;
        1692: s4_angle <= 25;
        1693: s4_angle <= 25;
        1694: s4_angle <= 26;
        1695: s4_angle <= 26;
        1696: s4_angle <= 26;
        1697: s4_angle <= 27;
        1698: s4_angle <= 27;
        1699: s4_angle <= 28;
        1700: s4_angle <= 28;
        1701: s4_angle <= 29;
        1702: s4_angle <= 29;
        1703: s4_angle <= 29;
        1704: s4_angle <= 30;
        1705: s4_angle <= 30;
        1706: s4_angle <= 31;
        1707: s4_angle <= 31;
        1708: s4_angle <= 31;
        1709: s4_angle <= 31;
        1710: s4_angle <= 0;
        1711: s4_angle <= 1;
        1712: s4_angle <= 1;
        1713: s4_angle <= 2;
        1714: s4_angle <= 3;
        1715: s4_angle <= 3;
        1716: s4_angle <= 4;
        1717: s4_angle <= 5;
        1718: s4_angle <= 5;
        1719: s4_angle <= 6;
        1720: s4_angle <= 7;
        1721: s4_angle <= 8;
        1722: s4_angle <= 8;
        1723: s4_angle <= 9;
        1724: s4_angle <= 9;
        1725: s4_angle <= 10;
        1726: s4_angle <= 11;
        1727: s4_angle <= 11;
        1728: s4_angle <= 12;
        1729: s4_angle <= 13;
        1730: s4_angle <= 13;
        1731: s4_angle <= 14;
        1732: s4_angle <= 15;
        1733: s4_angle <= 15;
        1734: s4_angle <= 16;
        1735: s4_angle <= 16;
        1736: s4_angle <= 17;
        1737: s4_angle <= 17;
        1738: s4_angle <= 18;
        1739: s4_angle <= 19;
        1740: s4_angle <= 19;
        1741: s4_angle <= 20;
        1742: s4_angle <= 20;
        1743: s4_angle <= 21;
        1744: s4_angle <= 21;
        1745: s4_angle <= 22;
        1746: s4_angle <= 22;
        1747: s4_angle <= 23;
        1748: s4_angle <= 23;
        1749: s4_angle <= 24;
        1750: s4_angle <= 24;
        1751: s4_angle <= 25;
        1752: s4_angle <= 25;
        1753: s4_angle <= 26;
        1754: s4_angle <= 26;
        1755: s4_angle <= 27;
        1756: s4_angle <= 27;
        1757: s4_angle <= 27;
        1758: s4_angle <= 28;
        1759: s4_angle <= 28;
        1760: s4_angle <= 29;
        1761: s4_angle <= 29;
        1762: s4_angle <= 29;
        1763: s4_angle <= 30;
        1764: s4_angle <= 30;
        1765: s4_angle <= 31;
        1766: s4_angle <= 31;
        1767: s4_angle <= 31;
        1768: s4_angle <= 31;
        1769: s4_angle <= 0;
        1770: s4_angle <= 1;
        1771: s4_angle <= 1;
        1772: s4_angle <= 2;
        1773: s4_angle <= 3;
        1774: s4_angle <= 3;
        1775: s4_angle <= 4;
        1776: s4_angle <= 5;
        1777: s4_angle <= 5;
        1778: s4_angle <= 6;
        1779: s4_angle <= 7;
        1780: s4_angle <= 7;
        1781: s4_angle <= 8;
        1782: s4_angle <= 9;
        1783: s4_angle <= 9;
        1784: s4_angle <= 10;
        1785: s4_angle <= 11;
        1786: s4_angle <= 11;
        1787: s4_angle <= 12;
        1788: s4_angle <= 12;
        1789: s4_angle <= 13;
        1790: s4_angle <= 14;
        1791: s4_angle <= 14;
        1792: s4_angle <= 15;
        1793: s4_angle <= 16;
        1794: s4_angle <= 16;
        1795: s4_angle <= 17;
        1796: s4_angle <= 17;
        1797: s4_angle <= 18;
        1798: s4_angle <= 18;
        1799: s4_angle <= 19;
        1800: s4_angle <= 19;
        1801: s4_angle <= 20;
        1802: s4_angle <= 20;
        1803: s4_angle <= 21;
        1804: s4_angle <= 22;
        1805: s4_angle <= 22;
        1806: s4_angle <= 23;
        1807: s4_angle <= 23;
        1808: s4_angle <= 23;
        1809: s4_angle <= 24;
        1810: s4_angle <= 24;
        1811: s4_angle <= 25;
        1812: s4_angle <= 25;
        1813: s4_angle <= 26;
        1814: s4_angle <= 26;
        1815: s4_angle <= 27;
        1816: s4_angle <= 27;
        1817: s4_angle <= 27;
        1818: s4_angle <= 28;
        1819: s4_angle <= 28;
        1820: s4_angle <= 29;
        1821: s4_angle <= 29;
        1822: s4_angle <= 29;
        1823: s4_angle <= 30;
        1824: s4_angle <= 30;
        1825: s4_angle <= 31;
        1826: s4_angle <= 31;
        1827: s4_angle <= 31;
        1828: s4_angle <= 31;
        1829: s4_angle <= 0;
        1830: s4_angle <= 1;
        1831: s4_angle <= 1;
        1832: s4_angle <= 2;
        1833: s4_angle <= 3;
        1834: s4_angle <= 3;
        1835: s4_angle <= 4;
        1836: s4_angle <= 5;
        1837: s4_angle <= 5;
        1838: s4_angle <= 6;
        1839: s4_angle <= 7;
        1840: s4_angle <= 7;
        1841: s4_angle <= 8;
        1842: s4_angle <= 9;
        1843: s4_angle <= 9;
        1844: s4_angle <= 10;
        1845: s4_angle <= 10;
        1846: s4_angle <= 11;
        1847: s4_angle <= 12;
        1848: s4_angle <= 12;
        1849: s4_angle <= 13;
        1850: s4_angle <= 14;
        1851: s4_angle <= 14;
        1852: s4_angle <= 15;
        1853: s4_angle <= 15;
        1854: s4_angle <= 16;
        1855: s4_angle <= 16;
        1856: s4_angle <= 17;
        1857: s4_angle <= 18;
        1858: s4_angle <= 18;
        1859: s4_angle <= 19;
        1860: s4_angle <= 19;
        1861: s4_angle <= 20;
        1862: s4_angle <= 20;
        1863: s4_angle <= 21;
        1864: s4_angle <= 21;
        1865: s4_angle <= 22;
        1866: s4_angle <= 22;
        1867: s4_angle <= 23;
        1868: s4_angle <= 23;
        1869: s4_angle <= 24;
        1870: s4_angle <= 24;
        1871: s4_angle <= 25;
        1872: s4_angle <= 25;
        1873: s4_angle <= 25;
        1874: s4_angle <= 26;
        1875: s4_angle <= 26;
        1876: s4_angle <= 27;
        1877: s4_angle <= 27;
        1878: s4_angle <= 28;
        1879: s4_angle <= 28;
        1880: s4_angle <= 28;
        1881: s4_angle <= 29;
        1882: s4_angle <= 29;
        1883: s4_angle <= 30;
        1884: s4_angle <= 30;
        1885: s4_angle <= 30;
        1886: s4_angle <= 31;
        1887: s4_angle <= 31;
        1888: s4_angle <= 31;
        1889: s4_angle <= 31;
        1890: s4_angle <= 0;
        1891: s4_angle <= 1;
        1892: s4_angle <= 1;
        1893: s4_angle <= 2;
        1894: s4_angle <= 3;
        1895: s4_angle <= 3;
        1896: s4_angle <= 4;
        1897: s4_angle <= 5;
        1898: s4_angle <= 5;
        1899: s4_angle <= 6;
        1900: s4_angle <= 7;
        1901: s4_angle <= 7;
        1902: s4_angle <= 8;
        1903: s4_angle <= 8;
        1904: s4_angle <= 9;
        1905: s4_angle <= 10;
        1906: s4_angle <= 10;
        1907: s4_angle <= 11;
        1908: s4_angle <= 12;
        1909: s4_angle <= 12;
        1910: s4_angle <= 13;
        1911: s4_angle <= 13;
        1912: s4_angle <= 14;
        1913: s4_angle <= 14;
        1914: s4_angle <= 15;
        1915: s4_angle <= 16;
        1916: s4_angle <= 16;
        1917: s4_angle <= 17;
        1918: s4_angle <= 17;
        1919: s4_angle <= 18;
        1920: s4_angle <= 18;
        1921: s4_angle <= 19;
        1922: s4_angle <= 19;
        1923: s4_angle <= 20;
        1924: s4_angle <= 20;
        1925: s4_angle <= 21;
        1926: s4_angle <= 21;
        1927: s4_angle <= 22;
        1928: s4_angle <= 22;
        1929: s4_angle <= 23;
        1930: s4_angle <= 23;
        1931: s4_angle <= 24;
        1932: s4_angle <= 24;
        1933: s4_angle <= 25;
        1934: s4_angle <= 25;
        1935: s4_angle <= 26;
        1936: s4_angle <= 26;
        1937: s4_angle <= 26;
        1938: s4_angle <= 27;
        1939: s4_angle <= 27;
        1940: s4_angle <= 28;
        1941: s4_angle <= 28;
        1942: s4_angle <= 28;
        1943: s4_angle <= 29;
        1944: s4_angle <= 29;
        1945: s4_angle <= 30;
        1946: s4_angle <= 30;
        1947: s4_angle <= 30;
        1948: s4_angle <= 31;
        1949: s4_angle <= 31;
        1950: s4_angle <= 31;
        1951: s4_angle <= 31;
        1952: s4_angle <= 0;
        1953: s4_angle <= 1;
        1954: s4_angle <= 1;
        1955: s4_angle <= 2;
        1956: s4_angle <= 3;
        1957: s4_angle <= 3;
        1958: s4_angle <= 4;
        1959: s4_angle <= 5;
        1960: s4_angle <= 5;
        1961: s4_angle <= 6;
        1962: s4_angle <= 6;
        1963: s4_angle <= 7;
        1964: s4_angle <= 8;
        1965: s4_angle <= 8;
        1966: s4_angle <= 9;
        1967: s4_angle <= 10;
        1968: s4_angle <= 10;
        1969: s4_angle <= 11;
        1970: s4_angle <= 11;
        1971: s4_angle <= 12;
        1972: s4_angle <= 13;
        1973: s4_angle <= 13;
        1974: s4_angle <= 14;
        1975: s4_angle <= 14;
        1976: s4_angle <= 15;
        1977: s4_angle <= 15;
        1978: s4_angle <= 16;
        1979: s4_angle <= 16;
        1980: s4_angle <= 17;
        1981: s4_angle <= 18;
        1982: s4_angle <= 18;
        1983: s4_angle <= 19;
        1984: s4_angle <= 19;
        1985: s4_angle <= 20;
        1986: s4_angle <= 20;
        1987: s4_angle <= 21;
        1988: s4_angle <= 21;
        1989: s4_angle <= 22;
        1990: s4_angle <= 22;
        1991: s4_angle <= 23;
        1992: s4_angle <= 23;
        1993: s4_angle <= 24;
        1994: s4_angle <= 24;
        1995: s4_angle <= 24;
        1996: s4_angle <= 25;
        1997: s4_angle <= 25;
        1998: s4_angle <= 26;
        1999: s4_angle <= 26;
        2000: s4_angle <= 27;
        2001: s4_angle <= 27;
        2002: s4_angle <= 27;
        2003: s4_angle <= 28;
        2004: s4_angle <= 28;
        2005: s4_angle <= 28;
        2006: s4_angle <= 29;
        2007: s4_angle <= 29;
        2008: s4_angle <= 30;
        2009: s4_angle <= 30;
        2010: s4_angle <= 30;
        2011: s4_angle <= 31;
        2012: s4_angle <= 31;
        2013: s4_angle <= 31;
        2014: s4_angle <= 31;
	default: s4_angle <= 0;
      endcase
   end

   // [stage 5] generates a result
   wire [7:0] s5_res_1, s5_res_2, s5_res_3, s5_res_4, s5_res_5;
   assign s5_res_1 = s4_match  ? 32 : s4_angle;
   assign s5_res_2 = s4_swap   ? 64 - s5_res_1 : s5_res_1;
   assign s5_res_3 = s4_x_zero ? 0 : s4_y_zero ? 64 : s5_res_2;
   assign s5_res_4 = s4_y_neg  ? 128 - s5_res_3 : s5_res_3;
   assign s5_res_5 = s4_x_neg  ? 256 - s5_res_4 : s5_res_4;
   always @(posedge clock) begin
      out_val <= s5_res_5;
   end
   
   // functions ---------------------------------------------------------------
   function [7:0] absolute;
      input signed [8:0] value;
      begin
	 absolute = (value >= 0) ? value : -value;
      end
   endfunction
   
endmodule
`default_nettype wire

