//-----------------------------------------------------------------------------
// <simple_lsd>
//  - Simplified Line Segment Detector
//-----------------------------------------------------------------------------
// Version 1.07 (Nov. 12, 2019)
//  - Renamed the parameters <TAU>, <RHO>, and <MIN_LEN> to
//    <ANGLE_THRES>, <GRAD_THRES>, and <LENGTH_THRES> for clarity
//  - Changed the parameters shown above from local parameters to 
//    parameters which can be specified by a parent module
//  - Added automatic parameter tuning to avoid overutilization of
//    the line candidate RAM. If the utilization ratio exceeds 90%,
//    <GRAD_THRES> is incremented by <TUNING_STEP> every frame
//-----------------------------------------------------------------------------
// (C) 2019 Taito Manabe. All rights reserved.
//-----------------------------------------------------------------------------
`default_nettype none
`timescale 1ns/1ns

module simple_lsd
  #( parameter integer BIT_WIDTH    = 8,
     parameter integer IMAGE_HEIGHT = -1,
     parameter integer IMAGE_WIDTH  = -1,
     parameter integer FRAME_HEIGHT = -1,
     parameter integer FRAME_WIDTH  = -1,
     parameter integer ANGLE_THRES  = 16,   // (tau) max. angle difference
     parameter integer GRAD_THRES   = 655,  // (rho) min. grad. magnitude ** 2
     parameter integer LENGTH_THRES = 64,   // min. length of lines ** 2
     parameter integer RAM_SIZE     = 4096)
   ( clock, n_rst, in_y, in_vcnt, in_hcnt, out_flag, out_valid, 
     out_start_v, out_start_h, out_end_v, out_end_h, out_angle );

   // local parameters --------------------------------------------------------
   localparam integer ANGLE_BITW   = 8;   // currently, only 8 is supported
   localparam integer START_VCNT   = 0;
   localparam integer TUNING_STEP  = 16;
   localparam integer ATAN_LATENCY = 5;

   // following parameters are calculated automatically -----------------------
   localparam integer OVER_THRES   = (RAM_SIZE * 9) / 10;
   localparam integer H_BITW       = log2(FRAME_WIDTH);
   localparam integer V_BITW       = log2(FRAME_HEIGHT);
   localparam integer ADDR_BITW    = log2(RAM_SIZE);
   localparam integer COUNT_BITW   = log2(IMAGE_WIDTH  * IMAGE_HEIGHT);
   localparam integer DIST_BITW    = log2(IMAGE_WIDTH  * IMAGE_WIDTH +
					  IMAGE_HEIGHT * IMAGE_HEIGHT);
   localparam integer WORD_SIZE    
		      = 1 + DIST_BITW + (V_BITW + H_BITW + ANGLE_BITW) * 2;

   // inputs / outputs --------------------------------------------------------
   input wire 	                clock, n_rst;
   input wire [BIT_WIDTH-1:0] 	in_y;
   input wire [V_BITW-1:0] 	in_vcnt;
   input wire [H_BITW-1:0] 	in_hcnt;
   output reg 			out_flag,    out_valid;
   output reg [V_BITW-1:0] 	out_start_v, out_end_v;
   output reg [H_BITW-1:0] 	out_start_h, out_end_h;
   output reg [ANGLE_BITW-1:0] 	out_angle;

   // applies Gaussian blur ---------------------------------------------------
   wire [BIT_WIDTH-1:0]       gau_pixel;
   wire [V_BITW-1:0] 	      gau_vcnt;
   wire [H_BITW-1:0] 	      gau_hcnt;
   gaussian
     #( .BIT_WIDTH(BIT_WIDTH), 
	.IMAGE_HEIGHT(IMAGE_HEIGHT), .IMAGE_WIDTH(IMAGE_WIDTH),
	.FRAME_HEIGHT(FRAME_HEIGHT), .FRAME_WIDTH(FRAME_WIDTH) )
   gau_0
     (  .clock(clock),         .n_rst(n_rst), 
	.in_pixel(in_y),       .in_vcnt(in_vcnt),   .in_hcnt(in_hcnt),
	.out_pixel(gau_pixel), .out_vcnt(gau_vcnt), .out_hcnt(gau_hcnt));

   // 2x2 window --------------------------------------------------------------
   wire [BIT_WIDTH-1:0]       stp_patch[0:1][0:1];
   wire [V_BITW-1:0] 	      stp_vcnt;
   wire [H_BITW-1:0] 	      stp_hcnt;
   stream_patch
     #( .BIT_WIDTH(BIT_WIDTH), 
	.IMAGE_HEIGHT(IMAGE_HEIGHT), .IMAGE_WIDTH(IMAGE_WIDTH),
	.FRAME_HEIGHT(FRAME_HEIGHT), .FRAME_WIDTH(FRAME_WIDTH),
	.PATCH_HEIGHT(2), .PATCH_WIDTH(2), .CENTER_V(0), .CENTER_H(0) )
   stp_0
     (  .clock(clock),         .n_rst(n_rst), 
	.in_pixel(gau_pixel),  .in_vcnt(gau_vcnt),  .in_hcnt(gau_hcnt),
	.out_patch({stp_patch[0][0], stp_patch[0][1], 
		    stp_patch[1][0], stp_patch[1][1]}),
	.out_vcnt(stp_vcnt),   .out_hcnt(stp_hcnt) );

   // applies 2x2 differential filters ----------------------------------------
   reg signed [BIT_WIDTH:0]   gx, gy;
   always @(posedge clock) begin
      gx <= $signed(({2'b0, stp_patch[0][1]} + stp_patch[1][1]) -
		    ({2'b0, stp_patch[0][0]} + stp_patch[1][0])) >>> 1;
      gy <= $signed(({2'b0, stp_patch[1][0]} + stp_patch[1][1]) -
		    ({2'b0, stp_patch[0][0]} + stp_patch[0][1])) >>> 1;
   end
   
   // calculates gradient -----------------------------------------------------
   localparam [BIT_WIDTH-1:0] EXPAND = 0;
   reg [BIT_WIDTH*2:0]        gx2, gy2;
   wire 		      grd_valid;
   wire [ANGLE_BITW-1:0]      grd_angle;
   wire [V_BITW-1:0] 	      grd_vcnt;
   wire [H_BITW-1:0] 	      grd_hcnt;
   reg [BIT_WIDTH*2:0] 	      grd_thres_offset;
   
   // norm check
   always @(posedge clock) begin
      gx2 <= ($signed({gx, EXPAND}) >>> BIT_WIDTH) * gx;
      gy2 <= ($signed({gy, EXPAND}) >>> BIT_WIDTH) * gy;
   end
   delay
     #( .BIT_WIDTH(1), .LATENCY(ATAN_LATENCY - 1) )
   dly_norm
     (  .clock(clock), .n_rst(n_rst), .out_data(grd_valid),
	.in_data(((gx2 + gy2) >= (GRAD_THRES + grd_thres_offset))) );

   // arctangent
   arctan_calc 
   atan_0
     (  .clock(clock), .in_x1(gx[BIT_WIDTH -:9]), .in_x2(gy[BIT_WIDTH -:9]), 
	.out_val(grd_angle[ANGLE_BITW-1 -:8]) );
   
   // coordinate adjustment
   coord_adjuster
     #( .FRAME_HEIGHT(FRAME_HEIGHT), .FRAME_WIDTH(FRAME_WIDTH), 
	.LATENCY(ATAN_LATENCY + 1))
   cda_0
     (  .clock(clock), .in_vcnt(stp_vcnt), .in_hcnt(stp_hcnt),
	.out_vcnt(grd_vcnt), .out_hcnt(grd_hcnt) );
   
   // stream_patch for valid flag and angle -----------------------------------
   wire [V_BITW-1:0]         vcnt;
   wire [H_BITW-1:0] 	     hcnt;
   wire 		     valid[0:2][0:3];
   wire [ANGLE_BITW-1:0]     angle[0:2][0:3];
   
   stream_patch
     #( .BIT_WIDTH(1 + ANGLE_BITW), 
	.IMAGE_HEIGHT(IMAGE_HEIGHT), .IMAGE_WIDTH(IMAGE_WIDTH),
	.FRAME_HEIGHT(FRAME_HEIGHT), .FRAME_WIDTH(FRAME_WIDTH),
	.PATCH_HEIGHT(3), .PATCH_WIDTH(4), .CENTER_V(1), .CENTER_H(1),
	.PADDING(0) )
   stp_1
     (  .clock(clock), .n_rst(n_rst), .in_pixel({grd_valid, grd_angle}),
	.in_vcnt(grd_vcnt), .in_hcnt(grd_hcnt),
	.out_patch({valid[0][0], angle[0][0], valid[0][1], angle[0][1],
		    valid[0][2], angle[0][2], valid[0][3], angle[0][3],
		    valid[1][0], angle[1][0], valid[1][1], angle[1][1], 
		    valid[1][2], angle[1][2], valid[1][3], angle[1][3],
		    valid[2][0], angle[2][0], valid[2][1], angle[2][1], 
		    valid[2][2], angle[2][2], valid[2][3], angle[2][3]}),
	.out_vcnt(vcnt),    .out_hcnt(hcnt) );

   // common registers / wires ------------------------------------------------
   // state and output
   reg [1:0] 		     state;
   reg 			     overused;

   reg [ADDR_BITW-1:0] 	     read_id;
   // segment parameters
   reg 			     tracing, last;
   reg signed [ADDR_BITW:0]  seg_id;
   reg [DIST_BITW-1:0] 	     max_dist;
   reg [V_BITW-1:0] 	     end_1_v, end_2_v;
   reg [H_BITW-1:0] 	     end_1_h, end_2_h;
   reg [ANGLE_BITW-1:0]      angle_1, angle_2;
   reg [ADDR_BITW:0] 	     seg_num;
   // FIFO / RAM
   wire signed [ADDR_BITW:0] prev_id_out;
   reg 			     ram_wr_en;
   reg [ADDR_BITW-1:0] 	     ram_wr_addr;
   reg [WORD_SIZE-1:0] 	     ram_wr_data;
   wire [WORD_SIZE-1:0]      ram_rd_data;
   
   // state and data output control -------------------------------------------
   always @(posedge clock) begin
      if(!n_rst) begin
	 state <= 2;
      end
      else if(state == 0) begin   // search
	 if(vcnt == IMAGE_HEIGHT - 1 && hcnt == FRAME_WIDTH - 1) begin
	    state <= 1;
	    read_id <= 0;
	 end
      end
      else if(state == 1) begin   // output
	 if(read_id == seg_num)
	   state <= 2;
	 read_id <= read_id + 1;
      end
      else if(state == 2) begin   // wait
	 if((vcnt == (START_VCNT == 0 ? FRAME_HEIGHT - 1 : START_VCNT - 1)) &&
	    (hcnt == FRAME_WIDTH - 1)) begin
	    state <= 0;
	 end
      end
   end
     
   // tracing (termination) ---------------------------------------------------
   wire 		     cond_term_trace, cond_save_seg;   
   wire [ANGLE_BITW-1:0]     res_la1, res_la2;
   wire [DIST_BITW-1:0]      res_d1,  res_d2,  res_max_dist;
   wire [V_BITW-1:0] 	     res_end_1_v, res_end_2_v;
   wire [H_BITW-1:0] 	     res_end_1_h, res_end_2_h;
   wire 		     res_cond_1,  res_cond_2;   
   // condition
   assign cond_term_trace 
     = tracing && ((hcnt == IMAGE_WIDTH) || !valid[1][1] ||
		   (angle_diff(res_la1, res_la2) >= 2 * ANGLE_THRES));
   assign cond_save_seg   
     = cond_term_trace && (!last || (res_max_dist >= LENGTH_THRES));
   // update
   assign {res_la1, res_la2} 
     = update_range(angle_1, angle_2, angle[1][1]);
   assign res_d1     = calc_dist2(end_1_v, end_1_h, vcnt, hcnt - 1);
   assign res_d2     = calc_dist2(end_2_v, end_2_h, vcnt, hcnt - 1);
   assign res_cond_1 = (res_d1 >= res_d2) && (res_d1 > max_dist);
   assign res_cond_2 = (res_d2  > res_d1) && (res_d2 > max_dist);
   assign {res_end_2_v, res_end_2_h}
     = res_cond_1 ? {vcnt, hcnt - 1'b1} : {end_2_v, end_2_h};
   assign {res_end_1_v, res_end_1_h} 
     = (!res_cond_1 && res_cond_2) ? {vcnt, hcnt - 1'b1} : {end_1_v, end_1_h};
   assign res_max_dist
     = res_cond_1 ? res_d1 : res_cond_2 ? res_d2 : max_dist;
   
   // tracing (initialization / in-line update) -------------------------------
   wire [ANGLE_BITW-1:0]     up1_angle_1, up1_angle_2;
   wire [DIST_BITW-1:0]      up1_max_dist;
   wire [V_BITW-1:0] 	     up1_end_1_v, up1_end_2_v;
   wire [H_BITW-1:0] 	     up1_end_1_h, up1_end_2_h;
   wire signed [ADDR_BITW:0] up1_seg_id;
   wire 		     up1_last;

   assign up1_angle_1  = tracing ? res_la1 : angle[1][1];
   assign up1_angle_2  = tracing ? res_la2 : angle[1][1];
   assign up1_max_dist = tracing ? max_dist : 0;
   assign {up1_end_1_v, up1_end_1_h}
     = tracing ? {end_1_v, end_1_h} : {vcnt, hcnt};
   assign {up1_end_2_v, up1_end_2_h}
     = tracing ? {end_2_v, end_2_h} : {vcnt, hcnt};
   assign up1_seg_id   = tracing ? seg_id : seg_num;
   assign up1_last     = tracing ? last : 1;
   
   // tracing (searches for candidates in the previous line) ------------------
   // segment IDs of pixels in the previous line
   reg signed [ADDR_BITW:0]  prev_id[0:2];
   always @(posedge clock) begin
      prev_id[2] <= prev_id_out;
      prev_id[1] <= prev_id[2];
      prev_id[0] <= prev_id[1];
   end
   // selects the ID to be read from RAM
   wire signed [ADDR_BITW:0] pid_tmp;
   reg signed [ADDR_BITW:0]  pid;
   reg 			     found;
   assign pid_tmp 
     = ((prev_id[0] != -1) && (hcnt != FRAME_WIDTH - 1) && 
	(angle_diff(angle[0][1], angle[1][2]) < ANGLE_THRES)) ? prev_id[0] :
       ((prev_id[1] != -1) && 
	(angle_diff(angle[0][2], angle[1][2]) < ANGLE_THRES)) ? prev_id[1] :
       ((prev_id[2] != -1) && (hcnt != IMAGE_WIDTH - 2) && 
	(angle_diff(angle[0][3], angle[1][2]) < ANGLE_THRES)) ? prev_id[2] : -1;
   always @(posedge clock) begin
      pid   <= pid_tmp;
      found <= (pid_tmp != -1) && (vcnt > 0);
   end

   // tracing (obtains parameters of the candidate region) --------------------
   wire 		     pexist;
   wire [DIST_BITW-1:0]      pmd;
   wire [V_BITW-1:0] 	     pe1_v, pe2_v;
   wire [H_BITW-1:0] 	     pe1_h, pe2_h;
   wire [ANGLE_BITW-1:0]     pa1, pa2;   
   assign {pexist, pmd, pe1_v, pe1_h, pe2_v, pe2_h, pa1, pa2}
     = (ram_wr_en && (ram_wr_addr == pid)) ? ram_wr_data : ram_rd_data;

   // tracing (merges the candidate region into the current one) --------------
   // temp
   wire 		     cond_do_trace,   cond_merge;   
   wire [DIST_BITW-1:0]      up2_d[0:3], up2_max_d;
   wire [ANGLE_BITW-1:0]     up2_angle_1_tmp1, up2_angle_2_tmp1;
   wire [ANGLE_BITW-1:0]     up2_angle_1_tmp2, up2_angle_2_tmp2;
   wire [1:0] 		     up2_argmax;
   wire [V_BITW-1:0] 	     up2_max_e1_v, up2_max_e2_v;
   wire [H_BITW-1:0] 	     up2_max_e1_h, up2_max_e2_h;
   // results
   wire [DIST_BITW-1:0]      up2_max_dist;
   wire [ANGLE_BITW-1:0]     up2_angle_1, up2_angle_2;
   wire [V_BITW-1:0] 	     up2_end_1_v, up2_end_2_v;
   wire [H_BITW-1:0] 	     up2_end_1_h, up2_end_2_h;
   wire signed [ADDR_BITW:0] up2_seg_id;
   // conditions
   assign cond_do_trace 
     = !cond_term_trace && (hcnt < IMAGE_WIDTH) && valid[1][1];
   assign cond_merge
     = cond_do_trace && found && pexist && 
       (angle_diff(up2_angle_1_tmp2, up2_angle_2_tmp2) < ANGLE_THRES * 2);   
   // checks whether a new angle range is within the tolerance
   assign {up2_angle_1_tmp1, up2_angle_2_tmp1} 
     = update_range(pa1, pa2, up1_angle_1);
   assign {up2_angle_1_tmp2, up2_angle_2_tmp2} 
     = update_range(up2_angle_1_tmp1, up2_angle_2_tmp1, up1_angle_2);
   assign {up2_angle_1, up2_angle_2} 
     = !cond_merge ? {up1_angle_1, up1_angle_2} :
       {up2_angle_1_tmp2, up2_angle_2_tmp2};
   // updates start/end positions
   assign up2_d[0] = calc_dist2(pe1_v, pe1_h, up1_end_1_v, up1_end_1_h);
   assign up2_d[1] = calc_dist2(pe1_v, pe1_h, up1_end_2_v, up1_end_2_h);
   assign up2_d[2] = calc_dist2(pe2_v, pe2_h, up1_end_1_v, up1_end_1_h);
   assign up2_d[3] = calc_dist2(pe2_v, pe2_h, up1_end_2_v, up1_end_2_h);
   assign {up2_argmax, up2_max_d} 
     = dist_argmax4(up2_d[0], up2_d[1], up2_d[2], up2_d[3]);
   assign {up2_max_e1_v, up2_max_e1_h}
     = (up2_argmax < 2) ? {pe1_v, pe1_h} : {pe2_v, pe2_h};
   assign {up2_max_e2_v, up2_max_e2_h}
     = (up2_argmax[0] == 0) ? {up1_end_1_v, up1_end_1_h} 
       : {up1_end_2_v, up1_end_2_h} ;
   assign {up2_max_dist, up2_end_1_v, up2_end_1_h, up2_end_2_v, up2_end_2_h}
     = (cond_merge && (up2_max_d > up1_max_dist) && (up2_max_d > pmd)) ?
       {up2_max_d, up2_max_e1_v, up2_max_e1_h, up2_max_e2_v, up2_max_e2_h} :
       (cond_merge && (up1_max_dist < pmd)) ?
       {pmd, pe1_v, pe1_h, pe2_v, pe2_h} :
       {up1_max_dist, up1_end_1_v, up1_end_1_h, up1_end_2_v, up1_end_2_h};
   // decides an ID for the current segment
   assign up2_seg_id 
     = (cond_merge && !tracing) ? pid : up1_seg_id;

   // tracing (checks if there are any candidates in the next line) -----------
   wire 		     up2_last;
   assign up2_last
     = (vcnt < IMAGE_HEIGHT - 1) &&
       ((valid[2][0] && (hcnt != 0) &&
	 (angle_diff(angle[2][0], angle[1][1]) < ANGLE_THRES)) ||
	(valid[2][1] && 
	 (angle_diff(angle[2][1], angle[1][1]) < ANGLE_THRES)) ||
	(valid[2][2] && (hcnt != IMAGE_WIDTH - 1) &&
	 (angle_diff(angle[2][2], angle[1][1]) < ANGLE_THRES))) ? 0 : up1_last;

   // updates parameters ------------------------------------------------------
   always @(posedge clock) begin
      if(!n_rst) begin
	 tracing <= 0;
      end
      else begin
	 {angle_1, angle_2} <= {up2_angle_1, up2_angle_2};
	 {end_1_v, end_1_h} <= {up2_end_1_v, up2_end_1_h};
	 {end_2_v, end_2_h} <= {up2_end_2_v, up2_end_2_h};
	 {max_dist, seg_id, last} <= {up2_max_dist, up2_seg_id, up2_last};
	 tracing <= cond_do_trace ? 1 : 0;
      end
   end   
   
   // delay for obtaining segment IDs in the previous line --------------------
   delay
     #( .BIT_WIDTH(log2(RAM_SIZE) + 1), .LATENCY(FRAME_WIDTH - 3) )
   dly_0
     (  .clock(clock), .n_rst(n_rst),
	.in_data(cond_do_trace ? up2_seg_id : -1), .out_data(prev_id_out) );
   
   // RAM for seg_list (segment list) RAM -------------------------------------
   ram_sc
     #( .WORD_SIZE(WORD_SIZE), .RAM_SIZE(RAM_SIZE) )
   ram_0
     (  .clock(clock),         .wr_en(ram_wr_en),
	.wr_addr(ram_wr_addr), .wr_data(ram_wr_data),
	.rd_addr((state == 0) ? pid_tmp[ADDR_BITW-1:0] : read_id), 
	.rd_data(ram_rd_data) );

   // RAM control
   always @(posedge clock) begin
      if(!n_rst) begin
	 {seg_num, ram_wr_en} <= 0;
      end
      else begin
	 // starts inputting a new frame	 
	 if((vcnt == (START_VCNT == 0 ? FRAME_HEIGHT - 1 : START_VCNT - 1))
	     && (hcnt == FRAME_WIDTH - 1) ) begin
	    seg_num   <= 0;
	 end
	 // stops tracing and writes the integrated line segment
	 else if(cond_save_seg) begin
	    ram_wr_en   <= (state == 0) ? 1 : 0;
	    ram_wr_addr <= seg_id;
	    ram_wr_data <= {1'b1, res_max_dist, res_end_1_v, res_end_1_h,
			    res_end_2_v, res_end_2_h, angle_1, angle_2};
	    seg_num     <= ((state == 0) && (seg_id == seg_num) &&
			    (seg_num != RAM_SIZE - 1)) ?
			   seg_num + 1 : seg_num;
	 end
	 // invalidation
	 else if(cond_merge && tracing && (up1_seg_id != pid)) begin
	    ram_wr_en   <= (state == 0) ? 1 : 0;
	    ram_wr_addr <= pid;
	    ram_wr_data <= 0;
	 end
	 else begin
	    ram_wr_en   <= 0;
	 end
      end
   end

   // automatic threshold control ---------------------------------------------
   always @(posedge clock) begin
      if(!n_rst) begin
	 {overused, grd_thres_offset} <= 0;
      end
      else begin
	 // starts inputting a new frame	 
	 if((vcnt == IMAGE_HEIGHT) && (hcnt == 0)) begin
	    if(overused)
	      grd_thres_offset <= grd_thres_offset + TUNING_STEP;
	    else if(TUNING_STEP <= grd_thres_offset)
	      grd_thres_offset <= grd_thres_offset - TUNING_STEP;
	    overused <= 0;
	 end
	 // stops tracing and writes the integrated line segment
	 else if(cond_save_seg) begin
	    if((state == 0) && (OVER_THRES < seg_id))
	      overused <= 1;
	 end
      end
   end   
   
   // output ------------------------------------------------------------------
   wire [ANGLE_BITW-1:0]     swp_ad, mid_angle;
   assign swp_ad = angle_diff(pa1, pa2);
   assign mid_angle
     = (pa1 + swp_ad == pa2) ? (pa1 + swp_ad / 2) : (pa2 + swp_ad / 2);
   
   always @(posedge clock) begin
      out_flag  <= (state == 1) && (read_id >= 1);
      out_valid <= (pmd >= LENGTH_THRES);
      if(((( 32 <= mid_angle) && ( mid_angle <  96)) && (pe1_v < pe2_v)) ||
	 ((( 96 <= mid_angle) && ( mid_angle < 160)) && (pe1_h < pe2_h)) ||
	 (((160 <= mid_angle) && ( mid_angle < 224)) && (pe1_v > pe2_v)) ||
	 (((  mid_angle < 32) || (224 <= mid_angle)) && (pe1_h > pe2_h)))
	{out_start_v, out_start_h, out_end_v, out_end_h}
	  <= {pe2_v, pe2_h, pe1_v, pe1_h};
      else
	{out_start_v, out_start_h, out_end_v, out_end_h}
	  <= {pe1_v, pe1_h, pe2_v, pe2_h};
      out_angle <= mid_angle;
   end
     
   // functions ---------------------------------------------------------------
   // calculates angle difference between a and b
   function [ANGLE_BITW-1:0] angle_diff;
      input [ANGLE_BITW-1:0] a, b;
      reg [ANGLE_BITW-1:0]   abs_diff;  // this is not a register
      begin
	 abs_diff   = (a > b) ? (a - b) : (b - a);
	 angle_diff = ({abs_diff, 1'b0} < (1 << ANGLE_BITW)) ?
		      abs_diff : (1 << ANGLE_BITW) - abs_diff;
      end
   endfunction

   // calculates the squared Euclid distance between (v1, h1) and (v2, h2)
   function [DIST_BITW-1:0] calc_dist2;
      input signed [DIST_BITW:0] v1, h1, v2, h2;
      begin
	 calc_dist2 = (v1 - v2) * (v1 - v2) + (h1 - h2) * (h1 - h2);
      end
   endfunction

   // updates angle range [angle_1, angle_2] depending on <new_angle>
   function [ANGLE_BITW*2-1:0] update_range;
      input [ANGLE_BITW-1:0] angle_1, angle_2, new_angle;
      reg [ANGLE_BITW-1:0]   seg_range, range_1, range_2;
      // these are not registers
      begin
	 seg_range = angle_diff(angle_1, angle_2);
	 range_1   = angle_diff(new_angle, angle_1);
	 range_2   = angle_diff(new_angle, angle_2);
	 if( (range_1 >= range_2) && (range_1  > seg_range) )
	   update_range = {angle_1, new_angle};
	 else if( (range_2 > range_1) && (range_2 > seg_range) )
	   update_range = {new_angle, angle_2};
	 else
	   update_range = {angle_1, angle_2};
      end
   endfunction

   function [2+DIST_BITW-1:0] dist_argmax4;
      input [DIST_BITW-1:0] d0, d1, d2, d3;
      reg 		    max_arg1, max_arg2; // | not registers
      reg [DIST_BITW-1:0]   max_val1, max_val2; // | 
      begin
	 max_arg1 = (d0 > d1) ? 0  : 1;
	 max_val1 = (d0 > d1) ? d0 : d1;
	 max_arg2 = (d2 > d3) ? 0  : 1;
	 max_val2 = (d2 > d3) ? d2 : d3;
	 dist_argmax4 = (max_val1 > max_val2) ? 
			{1'b0, max_arg1, max_val1} : {1'b1, max_arg2, max_val2};
      end
   endfunction
   
   function integer log2;
      input integer value;
      begin
     	 value = value - 1;
	 for(log2 = 0; value > 0; log2 = log2 + 1)
	   value = value >> 1;
      end
   endfunction
   
endmodule
`default_nettype wire
